��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!��Q�"u�b�c�#3�-{_sh�o�vAg~�r)�t~IV�z�������U��d�ф~����p�1!�΋;Dvn��I�?��]����W���' 㴟��Gn��:6�r���p��VL��*(o���6v3��'Ytp��:;�[���!P��~�|M*Ęj2�B�[�b�x�L(����A.����4��i�%�!�>����O�	
ߗk�J��I�z�]�c���x8��H��Z��{_��iЊW���5ºvB�s~,ptQ���}�L<v��e4�����3dJp��L�8H�@7��G���ږ�3xZVP�Xr�][�@���rah����f�����6�Lq�2,ߏt�Ĵϼ	���6�э�|�����B�3|}s珇�EH%ō���!�X��KȘG%�=p��SjT���O�vq�M�4�H��H�Ǉ&���M�6��v����
#U���:�Q�kv> ���mz�� |��/�Xh��:e[�#�մ�.B;O.��Oz���t ��c���x�6���v���?�֋d���=L���4_�?GQ�.��V��?oj�s�g�7���ϾU};ɀ`;�4���(~�MǓߥp$���"��dZ0o�v�T��^�v!��$0j?�s�����XI�a�f2�[���ٹ���م�uLꏯ<>x�2`�J�É�����d�x����e������k	����UvЅ��Q��j�`�ϋ��GmJ��ɼی(y�3�`�����x���B,'u���/8'�QL&�v��H��2���2�()Ȕ�7� �M��O ��� 1�+�44΄,�H'u$�5�=�7ȸ���<h�<�V�QK�}�Y>�K-85I��ޥ�9���b�j��}�d�܂��Y�kí��K��Gn�*TȷG١��3	[G;�\5�I���(����<��Q��V�ea���}ڌ�� ��1���d�O��{��nrm؊(�p�Y���U�m����]�cS�GN�f�U*�qMC�%`zh��g(>����;�Ӏ�sqS�I)ŢeD��8�>z��4%��짐��R%%F�%��짐�(�N���P�7H����>��E������y�.q�Q�Ҷ�dǙ��
��A|������7�ݒ}dZ0o�vʱ3������6��n��`���n=2�����(å
�A뫰v]uR���C(QGŎ·�K`������l<�Qudw��|@�M���5^s桃��k�Ĳh;�E{-�>�����B�ժ����J�A��\�${i���~�;�m^$��
�/��,�R_cb�
#2y��g??���CM��5�Sz��6�Lq����P/�[�CM��5�Sz֞��� ��� @����eGfFXջ�hʢ!�5�	�����ތsȸ�"rR��(�ٱ�W�I�z�]��&���V�g�TI���P��mgA��k\�����"�9i&�Q0�u���%��짐�(��v�r�]s�ES�T�<L�*-��pޒ�.��P]:�K!��]#5؝��Ү���<Mz�0�4��3�>=���#,J�l�/f#�}N9�h�{JB"���y�#=�h��M���5^s�=�kN�j�����ʂ�)Af@�k�&�厏�c���Z/2�sȸ�"rR�P�΃�F��t�Ძʃ���#_��⋬n��2%0���K+�,x�W��.��贅����c�Ѽ?���FCx��!�`�(i3}C��uo	�l+%��xC��=��:67�,���%�����	����o����ry�TG,���%����(��X> r[B1Y������Fz�<4f/J8�<}�L�Wa��Ĩ4�/T��ê�Kq���a�S�P��3,.x�Ȫ�>�B�HCڰ������c�H���ׇӭ��5�����}Y�e�E*'/	�7.����f��%
�������FP��cC�Ic9S��D�j���r��܊F`��j�.S2ׇӭ��I����d��r�b+ǯ3�4���G2���*�)���K����c�!z�i	'3�=٪	�Z�I�C�8%~��im��ғ�;ab95c�����m��!���"h��1���!im�Ia�|�����>ր 6���%k�����T�:�g??���9��xqw$FD��N�3��뙾�SYO�i�%��!�r����2��O�&cj=�׶�@�$Y�*#�IQ܋�9�2"�!�`�(i3C�A<�Z�̳P�ߙ[qwQ{>�붋"�M~O���ƻo2j�`$|�ku\ad����6�z�
^9�*�l9yt��g4sȸ�"rR��0�&�ͭ���<My�zk98�5��W(��ɗ�s�
>{J�^C���m��o30�@C7��G���ږ�3xZV���)n?����뺨����>=���#Y�J����x���Uͱ�YxM��}�!�`�(i3�Y��nkMM��m�7�TG�>{=�b]!	r��m�z��b6������P��y�#=�h��M���5^s�"��FlXz~�Gy�'W��	]�	���D��ܒ�����[m	���Ʉ �����#(L�̷v2�j!�`�(i3Y�Q3�tY�Dy�-����F>����٭M�3�9��)pZ���b�a�WX3�T?ې!p���.��Щv<�<��hK.���Fz�bˑn�9�Ƅ^�=�]�_Jz���j
a�I���;% ���WyffwA�!�`�(i3�"��kyB��ljrk���Q�4IS88��9/���`���6j��p����]n���Q�lH�K&�\�4�ʈKk�IkY�G�ׇӭ�ц�'T���+Y�������l5,/���=`�*嘌\k%��Ns�$���^O��<!�`�(i3:�8���V����
�?<��2������p����]n��؜v�4�oe��t-߱�~�jf&�~�7��o���̄1��7���Fz��V�52SG���Vd�'�K��{�!�9��&A�����˛q!�`�(i3�LQ&��w+K>�_��c����}��[�P5����N?4Y�1V*���p���h�n�ഛ�r��!�`�(i3:�8���V��yoZ�P/��B���- ��[T� c����}���R�-�촎LQ愥~�����8�/��y:����Fz��ݓ�W���Wtܓ��o5xM�����?��9)7�S�����f���;�[!�`�(i3�LQ&��w,V׋jŀ����Dg�D�M>b�B���Zb���6�z�
^Hj����85I��ޥm�>�
 !�`�(i3:�8���V��A�,�4���/,��YHiJU�4�B��ٴ���j>��	��x<�b�Kf�������1EZYq�A�G�+H�pVl�x�7~�8!��� �)cΝ���g??���CM��5�Sz��*^QP�o4�m�ρ�4��	���z�K�fC���4M=���^���Fz�2Y��kک�@ɤ��ӄ+����<�r<��ou���&�����Q�W0jD��D1��n	�I]��Q*7��0�c�k2�}�sȸ�"rRY�5c�P))�jf&�~�7���p�J�����qZ��B[��_Um-V|S��=�=����ly/Z�Ns�`�ϋ��Gr
6����8X�˞�DG!�`�(i3�N�����>��#����2��cF�a\Y������t潅�����c��R����<Fl�Ř#7⸠z�V[���KdyQ��G�T3$!�`�(i3\zgn�K���&�mN-�07����F��k.J���g�|R��qB$e���)\EH�a���\�����
�Z���R�t�r�B���J{��!�`�(i3q�\E��0\��M��ړ'�al��p�~����p|K�mb�Xm[ �tf�A�����KNJ����� O
Ү��p75傟������t_��?�T���� �� \���q���~����[T� ��~��Αu#��Ͳ0�nh1=2��j��Z&��Ûf��O�.��+Y�B�&�%b]���$��Q;�]�1T��v���_�G��Gq{�f��a��{oS���%�a�����v��C�Gx�-��;ۂ��IÙ=�H��A��@1�
Ү��p75傟������t_��?���͈vLG2A�����ofv\y݅�ebÆ����޷�ס\���|K�{ߝ�t&REϞ]t��):����:���M��A���va�{����}����Y�Q�ki���cj~GM���Hc�@!��^�x)1�d�X�VM�����a�"�_���˥óM�˄Nc�r5�М`�@~��6��2��{�&>�_���6N�����=tUF����VrG+���)Uk�:��3���ne66�v��G�x�c�f�,b���開p+���`N���:�_���.�\�:���M��_(����@N��B�)Y��|K�{ߝ�;ª�����Q�u���Ifp`��<�W�C%c�����<�W�C%��b�^��ȭ�n�h��� v#7�K�=I  ����vȭ�n�h��� v#7n����K�����"��y�LN��K��g����R�<�W�C%c�����<�W�C%����_Wr��;���EWr�L{1��ox ������ �i7�sp>��w��sT��;���EWr���G����IÙ=�H
,�L�FӉ�w7N]���Ο2�K����3S4Wi�Baz�Ҽ���y�]���m ��-C�8�w����L�w�wr�4�V���jF~���F�v�*�1-0b���B���kDw|A��>��y�䃶&f��p�|�q��r/��5Տ�E`���_��	��\��g�p>�yn
V~$L�
�k���۪	�}a+J���k�����3�}@
-��[ȴ� �0�|���|K�{ߝ�2v�6�) �YR�42������:���M��A���va�{����2��� ��b�FP&T�p�lq�zL͊�q��C���岎� �1x�it�3�,#C~X��WG �����n�O�V��'[��uj}��8�,�G@�yLx(�i��/R#��`*�pv�r���Su�����f#�>���0;�Se�W@�óM�˄Nc�r5�М`�@~��6��fn=b�#O!��&M����ቸC�g�vUC+
]/R����3P�d�8!��vp�P}��O��^��mi9�g#���)��(0�w7�'n�^0o�:M`��e���im�����O�m������uH/Q����F�)�o?��?�Ddh�hq�ǆQV�� �h0�Y��A&�����jP�k׏�����M����8�&����+�`|��߉���_��V��E��a��óM�˄NO�7��Kq�c��ē��ľ2�ʓ�d�X�VM�����a�"�'n�^0o՘W��.�r����m�q� ������ �i7�sp>�Z�	�і�F�2��SbR��*H/Q�����Lm�yPǆQV�� �h0�Y�T��2�k�׏�����M����8�&����+���"%�i�;+HV�x��C�MV���t��tZ��_��V�V��>�����3P�d�8!��vp�P}��O��^��mi9�g#���)��(0�w7�'n�^0o�:M`��e���im���9:S�-M�O��~��Z>H@��4���ޡYB�R���>_�Z>H@���X~�� �4�04�jf�9��o�����Pm�|��1�gU��VB�����2��~ȭ�n�h��� v#70=$��_��A�F�7���3�GXS����E@��~���($�J.���
�L�Xڈ*-�kЄ�0v�J�NIyH\90\d'8�6�Pr"?uK!�����
; ���Y����=�\ǁٲ"q�Z˻r���5傟�����̝�wz�҄`�����'p�@�5傟������t_��?�GN0���!t|Y�f�s���N�k ��{m{Q�'g��|����ķQ�xO�ȭ�n�h�>�(BΫ�yp��Jy�t���Hhqu!���5�Nn���4L"�+�va��2{a�t P��p�U��o.��:��F��CǍԽB��'n�^0o��Ϊܜ��8TJ�����[T�)���y���OJHn��z��r9�3�B0)5�6.�/'�����W�^ֻ����XP��Ȇ<�qp^S��j.Z��$�sӢ�]3�����c��(r$����G[���0N������Y��,aAx��[U���z-j>yR�_o��ӳ�Y�
��M�P�zL͊�q��G�D�� ��o݆g��Э[�}��|�Q�iӻ�����.u-j>yR�_o�$�R�n��5��8�t��\�v�[������ڰN�& ��݊B\���̠ӷ��k2(
�D�lnA:�H�b���:��k>��'�@�TLN��=�u���i�)_�hil�C�����/*8���KP�i�IÙ=�H=Ӕ��()�1��b�:���rw��)^G�<�zL͊�q��j�[���'�`Uv��*(l��(�~�������k��whil�C��v��NrY��'��	�'n�^0o��W���M����Оy�*(l��(�~�������k��wK�]�Zw9=Lٽ����H�br����q{�f��a�:&�>��sH�2Da���`�M7Э��'D��h\e��6ڿ ����5�P���q�ِ�W���~*.�P[k�KW�*�	S,�d;vt��^_�V-��&'�ɀxm�������x���hAJHn��z�_c)���8��t���i�Oa�b��~��钏b�n���\���e�Q;���gq�IÙ=�HԹ��X��`w�~ڽwKl9
ya�Q{�K�-k/ /�:y�0�6�]���~����_j���=���a����Wo��̗�����H��@Ő��t��[=U�Z硘�`�Jk�IT�f|��P�����ʜ耚ҵԼ�\�v�\ !�d2�j�����PJ���9�a��C����\ԥ���u��TH�i$1x<�`�Oķ{y(����5�'n�^0o.�g���D�T̻6��v���[�SӠ� �9g�M�G�nʏ�(Z�ϯD�x�&��?GQ�.�,��o��h�76AyW���j�bB����^_�V-��&'�ɀxml�4��H���FÖ<^�q{�f��a�1��]2<�	=T�"E&��� ���yoZ�P/�]=a}��:��e��q�탯;\߰��V���
4�B��ٴ��
Y���}�Zs��as��5�"�r�x×v�XȪ,@�&>�JHn��z���hU��9�OZ+L�ʜ%�j@c�X[�\��!?�d���&�m6
�DR����ʺ�?���5��tR�&@>$!�u�]aL�ɜ���F)��`��z � �o*�voj�N�)�\x�s]���uC#���3Y���� �i7�sp>�{ƕ��w��\���\ ����@�!I/���P�>һo�%�ˏ8[$0�����|w"�_%�C��~�&A��`�����i�t�<�<俇d(�D-rB}VGڝ��s��WC�B8���9&	;�RP$W��q�b��'n�^0o�+#�K>��{�TNJ?�s�E(��6�ג�Û�����6�z�
^��2��Q�-���!Z�M�I����&A��`�����i�t�<�<俇d(�D-rB}VGڝ��s��WC�]��T&�t��Y�I��q{�f��a�:&�>��sH�2Da���`�M7Э7l��A���;��|BT׺Ò�<W�,C%���=�*��g�Ҙ�%Z_0@>$!�u�]aL�ɜ���F)��`��z � �o*�vo��sK�+�R��-f�u;5B5Y+� �i7�sp>��>9UW?8����V���Zy�>�@�מ�u��Ϣ�͹sC�MP7�B�J���1��b�,�MGuvh:a�������-7 �3�V���C��\����V�D���Kb���=���aٚ�o����6��/�6���� 9�������z�Ba����	#���,�+V�RDFR7�Y����0r����
���E�/$z{�Ѿ��h��#���%��#i�~cG���l�4��H���F(�E���/ښ[TJHn��z���YG�s�p$C���<��3�
W��1&&����$j.����.��79=��)^>�b*b  �H�,3�V���C��s�wWIÙ=�H�&8���l�mq���)�:�:O����6#�|ސ�r+�\�(��q@���TL߷�q5�ˉ�Ĭ	4�������x�jk��=y�/�xg�T��-7 �3�V���C�Y�i��x4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5Ғ�>S�8�dy��{W(l�4��H���Nx�W�^�U� ���_#8��shƻ9��[�>�q�E#�UJ�#��Iam�D6�U6qW�'n-i�& ܵz��O's;o@�1�9���9M/��:M/������;#���,�+V�RDFR7����_�b狡����
:�
5���4�~wD[����#9Fy7GD@�F��q`E�cvR+G
WW�r>1�C�G��$���
G�|�!<��l�
Q:Õ�)X�J�$�R�n�&�ގ/[ ���=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wI^+������_�����kf���Jx�]�V�����TI��ԑ�g��@��C$����}��yoZ�P/�i;@��\q.�YF�L�U���;�A+b���5,/�C�
؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U��aVN�+�S��t��)k�-ohHeg��|����s�ݺᣄ��C�W#@-�ʳ87��Q7�j�!��>��&pR��a��\�}1�-7 �3�V���C1
&���4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5Ғ�>S�8�dy��{W(l�4��H���YM�z}�؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U�/��2��'���ߌ[R)Ms	[�����-�2�{�OF8w?pª\��3͗I�+O��P�mO��'��U'j��p�U��o.�14�~�Xo��X���d�٣��c�A�L'b-a��K�aU�uC��v��{�'p#I^R)4�����5�2D�3����hV�:��ڴ�IÙ=�H�&8�����f���V�RDFR7��_���׍)�L�m�M�j`�;�_�2��B�>KJ��|�d��ķQ�xO�����y�� ː��+�w��IQ]~���+�#��V�d����Ԛ�ނ{�!��H�q�&������a
��20��4�|75Ol`V)�l֐�?���q.�����'��Ӥ�nq�IÙ=�H(�Y����>��NJ/��!�#��W+Δ}M��R���q{�f��a�:&�>��s��l�
Q:�A�;#�tױ�1���v�;)����=���aw��@�G��o�������HX�r	�y�L�G�I�[U���z-j>yR�_oݧG �ŴP��CnUc?��d��\�v��wc�}�![=���[](U�C��z��
������y��ٓA�ln�~ �i7�sp>F@��uݧG �ŴP��Cn��Y0C8�}4];ˍH���]&�HF@��uݧG �ŴP��Cnլ���4�L�U���;��n�^-@��M�fIÙ=�H�&8���l�mq���)�:�:O����6#�|ސ�r+�\�(��q�����N�l��u@����-_:�?]#���,�+�B�M�5���&�>,L��]��rň�����r���aM"��N�߄�4�X�)Х��؊�K�H��\�vūx`��:�=���[](U�C��z��0�<��_MÕ�)X�J"��Q����%�8j�<1�9���9MȎ��Mƀ�~'��u��m�.��H�c��1�%�e��G�b�<��]5���\�v��:Y��z��Mm�����X���n�{܎�)�V�H���!n}y���q���U�6�£p�=^�?GQ�.��V��?ojʣ='Xhy����A@�č�Y���S�)37J*uc�A�L'�f?S��ӳ�Y�
�ߪ��wZ�n��[��{_8�Y��=�}�Vݨ�%�fĀ�[�}��|M�9W2�R�E$OK�/�k�IkY�G���VѿZ� f�Lu�ms|d_!�\�<��z��}�0z�cUL���gM�6��A+b��ü~���U��g��U-�ee�@Rv����my$�N��lثl�;c����Ew(�A{d�F��M�9W2�R�E$OK�/�,�	��E"��VѿZ�R���O�C;=B>�ǈ��\�B�ҋX������S8�����)�dB%���O-�#���[�� ��q�%a(􆿳�tP"7��%e��0�UX�Pp42JF�Z��ʝ�>	���n�sӠ�k-q뚸�d���A�Pf�d�:h}�"+�{z �g��\�F�s��M_����
�?<N�Y�N�rb<��z��}�<ͧ�:|C���m9�/����Ew(�9V(;�&���܀�fH�k��v�~������]�!��	Ǹ�y85�V�9cޅU��9؜�%��Wǖg3ȓ8���/�l|�*"k���(ӈ�����w����>��5u�Qkgw��.:� tN���&�%_�DO� �Q�c�,e(}�_3#ڸZ鎬����Ĺ#{���t���@�����%zsӠ�k-q�Wv�A��1=ƌ�F�Y��D�n҃���:'�_���wg�!n}y��p�VU��J}\�=��Ӽ��2��}n	�Z^�t���,2����X�kX������`4�E%v�~������]�!���\B��V��PV�)ڶ�|ceJ�z��eU�e�����T�2���%,J�l�/]��-5L�S|��)����\�6�(�_3#ڸZ鎬����Ĺ#{�������犃�8�Qt�z��eU�e��������Dg��y��tqӴ����s��8�M���e���96��`��Лv�~������]�!���\B��Vjn.����Ϙ�J|�Qz��eU�e��������Dg��y��tqӴ����s��W�u��ó}����w�q��N���OG��_3#ڸZ鎬����Ĺ#{��2A���ϻ$�Zkԑ�]�Jg����-c �ЄW:l�mq���)�:;o�������=VU�����WΓ�Y�mݶ���č�Y���S�)37J*u�,�JL�������d)N�UE�B*�2���u���d���=A�2�S|���f?��� <���eW��H��ě�5/U�rQ��3c/��!`����J��<��z��}�<ͧ�:|C���m9�/s9}B�Ź��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,������[GL�����K+I�\�q��N��f�;�>)�~�`�0��|��].��'���Xw�����C��Z_�� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j����H��[n��B��X���WΓ�e'��ǩ����l�u+�v�~������]�!���\B��V�e9O��g��$y�z��eU�e��������Dg��y��tqӴ����s��~�̳o�"�D<�4_�;��	��Z\�i�æu�Q_�}{KS�)37J*u�,�JL�������d͇ :�s��]�Jg����-c �ЄW:l�mq���)�:;o�����p�ǔ|�b�ei�5/U�rQ��3c/��!w=����^<��z��}�<ͧ�:|C���m9�/�!������ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����&�2 ���������x��lV��(C6	�YI܁���!n}y��p�VU��J}\�=���T�<�����Z1~�g]�I���B��&���a�%�j@c�}������[
]&M��j���$5�}�����q>�~I� �_3#ڸZ鎬����Ĺ#{���Wl
% ��)ʒ�"��/8'�G~+�3;��\���\ ����@���d}�80�[X�b\g�8>!��J�0N�
���	�Bz���tU`f�g_3#ڸZ鎬�������(���R2�sW��t_-Z��T�\ �͘�f��p�b�z'hۉ)s���Ħ�q��Z1~�g]�I���B�龈4��G	������t4z��w���*#�IQ܋[���,d�܉-`�6�����Up��^��0� �8k>6s����]�!��	Ǹ�y85���~�h�Sü~���U��g��U-�e?�:�Z%�~kE#z��eU�e��������Ӟj��s �׊�8²u�8���=ON��t*�[P{C�#^r�3P���WT�j
�I��w��,�9���������a;�/8'�L
�2�Ot�ky����R� -�*3fN&����6��Ҡ��Nx]<	���rѮ�7]�8k>6s����]�!��	Ǹ�y85�ӓ��������@	Q��"X��[���`m��O���U4��{2l���^���@�d�_C�VJ����̕���(��hG�U�Ƕ�2��c=�_R�0��=��d�����caEyF�8ơ�@IE�U����S8�����)�dl�4��H���t_-Z��T�\ ��Sv[J�1ť�}<�&�/8'�G~+�3;��\���\��k�zph5)�� ��լ���MR�Ӝ�n����։�s/�yf��nͼ<�TD��x��3�]�����_�sL�jGC��w3�Z.��	.�V�~�-�r�e�L�]�തJ��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����Hg8l�6o���m�D��%�r �&M��y��Iۯ�oR���7�m��=�Ғ"_��5&���#�{�0;�}8�yaô��
; ����`���ś���e�7��(�kp�f�-���	ڐ�� Y��R�5����`K�y �谝��X�e���V!���IÙ=�H�SA���4��ɥ����%�a�HL����rm��U}�	KݗZ:���'n�^0onɌ����n������ɥ����%�a���.����^hq��:�}0�st&���\�v���T�©@���U@���:��F�Τow��@�5����`K�8dn�����bū�R��_�}���\�v�Fp~�]���s�b�a��wq�,���Hb^�G��$~������͌4s+�ny�H�5�o��r�i�H�^ֻ����XP����U�5Ϝjw$��$�ɋ��ă�s��z~�;�8dn�����bū�R��n���,�,���ۭ(��~T���ٿ�n�P�������h=�NWy1IPt|Y�f�sB�i�y�\��\�۟�-?�d���&����{ԕ�h7�{`���@�	��h;E����Y~��`�J���]�=�JHn��z��T��e�:0���ͭqRmHX���׫�J��;5B5Y+� �i7�sp>F@��u@���U@���:��F�b��@�zL͊�q��MQß�òo�P2}�).;��L�O#t����n��]ߺ�`@ZWH]�+��G=X��[���J2~M�G�}�+����+u��)_�������h[�f;q�s;5B5Y+��2tCH����,=3���Z�����Oy�����k2(
�D�lnA:��2Y���g��v�x��� T2��zL͊�q��T��Db
�o݆g���V�RDFR7�z�k�Bm��y?h�g&2�(K��ӿ����
Ym�����俧:zvkZ���6�� ���S%�eL)�1��bMI�����^ֻ����XP������a��l)�1��b�:���rw��)^G�<�zL͊�q��j�[���'�`Uv��*(l��(�~�������k��wh0%���dҺt��J��#Y��Ѽ�\�v���'ٍ&�cx�T �SNÕ�*lSf�IO�Ÿ��t+���/��2��w�\	_S>�xH���B){a�N*��XP������<����Dg��y��tq����A��(o�FP�١�&Y��V�$�Ƣ�/몱z���ۀm{�+{*N,=����/�C�ټ�)_����q{�7��)��}�OV9�a��j=IÙ=�H�Z�f�-�i��м8jqY���SހS�ɋ��ă�s;�B�;5B5Y+� �i7�sp>X�X�'��m�Ȕ�1���c]���;�"�!1�U��`__��g��|���y�~��ۢ��9��i��^z\�{�TDHu@�w_���(8@���c]���;�P�����ʜ耚ҵԼ�\�vŠ�B��닶	��};J9��1@��
�b*���t��祣��G=X��1x<�`�Oķ{y(����5�'n�^0o�+#��D�T̻6��v���[�SӠ� �9g�M�G�nʏ�(Z�ϯD�x�&��?GQ�.�b��, �k��G=X��7Sx:��yi����S(���S~���)_�T��|�BE���`B�,�'`��zL͊�q��G�D�� ��|��vt۱���[U�˵�a��݌9�;����[�4-�By��R�i&�V����Sv� O`S�KW�*�	S��ڪ�����$�R�n�m.�>"�RX+�/�o�IÙ=�Hw?pª\��l�mq���)�:��j8HQ��e�z���V�RDFR7������`��I�t?�_��B�e�D�*�Y�p�Yч���Ҟ�+�����ڪ������,���-x×v�X�8����յ��\�v�]������_�sL�S|���f?��AJ��vNW�w��fD��o30�@C��iߗ�{�(s�O�+�t&p�10 @>$!�u�]aL�ɜ���F)��`��z ����cD��ʧI�8��_�$�R�n�a��X�F@�(����IÙ=�H�&8���l�mq���)�:��j8HQ��e�z���V�RDFR7��ᚌ��J��:sS89�*uT?�Х |�8�}7E��O��O
+@~`��)�j�����x�d���?��(�G�H����ܖȪ,@�&>�JHn��z���hU��9�OZ+L�ʜ%�j@c�X[�\��!?�d���&����L���Ȕ���U(��L�S��;Pc��W�w��fDkޖ��4\m��.��Cq֌B�4�mg[�X���sK�+�R��-f�u;5B5Y+� �i7�sp>��>9UW?8����V���Zy�>�@�מ�u��Ϣ�͹sC�MP7�B�J���1��b�,�MGuvh:a�{��<X��I^+������_�����������ĈL���U� ���_Y�B~�����sr���oJo�w���#�lT&A.����4mB�2�1��o�ʳ87��Q7�j�!��>��~�h/����'5��WPu/����Ӡ�w��2D�A"m�/��F����K��eqi�á[�6���l �����4��5���R3T�����N5@]0v㛿̷��\��yoZ�P/}�iw�VJ���C7��#"���FC� 4P/�WS��t��)g�ֆ�F���\�v�]������_�sL�S|���f?�Z䗵�wEW��(*���ǚ�-��P�0��)�!e��yoZ�P/Hx`Q����ʳ87��Q7�j�!��>���,z]-,��BpLÕ�)X�J�$�R�n�\�B-y\���=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wW�'n-i�& ܵz�?�o9P}71�9���9M/��:M/������;#���,�+V�RDFR7����_�b�W󛂀3��-7 �3�V���Cے̓&B4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5�A\���ޯL�U���;�A+b��Sa[����{؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U,��BpLÕ�)X�J�$�R�n�&�ގ/[ ���=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wW�'n-i�& ܵz��f�^q O1�9���9M/��:M/������;#���,�+V�RDFR7����_�b�W󛂀3��-7 �3�V���C�D��4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5�A\���ޯL�U���;�A+b��J��*��[J؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U,��BpLÕ�)X�J�$�R�n�+SR������=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wW�'n-i�& ܵz��~��&�g��|����s�ݺᣄ��C�W#@-�ʳ87��Q7�j�!��>��&pR��� ����"[�.(+��S�*���X:�*��ܟ^}4��q���Ab�%^��!��1�̷��\pRWl0E���n���7��/��2��'���ߌ[u��ND��]�!��	Ǹ�y85�>T
BFa@#>��  7h��� ��E3�]��a�����5�2D�3����hV�:��ڴ�IÙ=�H�&8�����f���V�RDFR7��_���׍)�n�,e�P���P����ӑ7�\�V�D���Kb���=���a��;O��+�	6?�.�
oُ���O�<�D���$Z;Ӥ�*!���5�Nn�>�lU��ti�4:$�a�� �ʨթnJ�D��n�,e�P���P���Pz�����������'n�^0o����y�]ެ\�+f$߈�vJVt�l�褻�sv���-q]IÙ=�H��D\	"�B a�޶�oo=S���?\��4];ˍH���]&�H�z%�ژ�(9�X��RS��uڜ3Jw6�
�Y���V���
s���?�������r���aM"��n�^���'n�^0o����SVc=���[](U�C��z��
������y��ٓA�ln�~ �i7�sp>5��aF�~B%���O-�#���[�ǋ舊k&�x�]�V����*�Yb}9k� b����;e5V�]C��m͡r��b  �H�,!ԱX�|�0��h�0��'n�^0o����y�]=���[](U�C��z����Ջ�/Cp�14�~�Xo��0���$��c����zL͊�q���19TH���m�.��H�c��1�A8���$����[�&�pR<�K�?d�����x�]�V���(c���^��?e�V0Z�m�.��H�c��1�%�e��G�b�<��]5���\�v��:Y��z����bH�H�"'�7�c�p&ĩ+Ã��Q�0�	�A�����<��z��}�צ:�)�]7�˺�9/���`���6j&���1D��ՁO�#dv�~������]�!��	Ǹ�y85�ӓ��������@	Q��"X��[����fbK7͍��|��W&":��^�o�AXҹvXI)63X����8��߇r�KӐ�9�V�d4Cm f�Lu�ms|d_!�\�<��z��}�0z�cUL���gM�6��A+b��ü~���U��g��U-�ee�@Rv����my$�N��lثl�;c����Ew(�A{d�F��M�9W2�R�E$OK�/�,�	��E";�����Jo�l�W��Q�@��߿�D����W�<��z��}�0z�cUL���gM�6�����;e5V�]C���\�Ķ��"X��[����fbK7͍��|��W&":>/�k�oc��/HG9�G�q*��$��J�P]Ĳ:�1�@ �~)�sQ�I��N}�}�����aK �|��].��'���Xw�����C�6�£p�=^V�RDFR7�m��p�0�f��ú"[Ʈ����{l�f|��rs�i��=29��a)�1��bMI�������"X��[����fbK7͍��|��W&":��^�o�A���A��(o�FP��XҹvXI)�F�Bm��^N��P�T<�t�S��{l�f|��:2QYeƈ �-u���k
?X!��RS��uڜ3A�g�ƨk��+ƣ��0Fo�!޳Nt�sVڌ����Bt��k�|��|��].��'���Xw�����C�;R�<kQ~w���~��ݏ1��𠛕!��L��KI�;�����Ig`i�ҋX����L$�����/�{��U��+�N"����y��,2�����^���@�c}-Wh�4�B��ٴ�F6_%v��w\�f@��<�Cr����Ig`i�ҋX����L$�����/�{��U��+8cR�F�㯆ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,�����Vt�%����"��#ߠR~36�{��B�ip��{l�f|��:2QYeƈ �-u���kS̅��|�B*�2���u���d���=A�2�S|���f?��� <�?W�&����t��!`(HYz�>�d�<��
�}����[v��{l�f|��:2QYeƈ �-u���k�����n� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j��a:��8<�I�3��
ip@55��;��CF�x&_3#ڸZ鎬����Ĺ#{�����U�^�"�� 1�	Q��,2�����^���@�d�_C�VJ����̕���(��h~���O��Q:���p�$�|��k<�<�`�hE���Mz��;��ҋX����L$�����/�{��U��+�����E)S��,2�����^���@�d�_C�VJ����̕���(��h��+��<ȫ� `�r��Y�Ȅ�f�;�>)�~�`�0��|��].��'���Xw�����C��Z_�� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j����H��[n��B��X���WΓ�BD{���p�պ����u�Q_�}{KS�)37J*u�,�JL�������d���J�l�]�Jg����-c �ЄW:l�mq���)�:;o�����G�̥}�ߘ����N�[վh��[�3c/��!?V#$~@!<��z��}�<ͧ�:|C���m9�/Ɨ@��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����&�2 �����&G|2-m�Y�Ȅ�f�;�>)��5�g��|��].��'���Xw�����C��*��z�)� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j��S��^1���k(�2��c=�_R�����t{�č�Y���S�)37J*u�,�JL�������d�`�%�]�]�Jg����-c �ЄW:l�mq���)�:�ۇT�0��e�zt�z��Al�q고�����f{ �$���{l�f|��:2QYeƈ �-u���ke�>��E۳B*�2���u���d���=A�2�S|���f?NԆ��-�ê�%�S��!���A���ՖC�͓Wԙ�"�F�%Q�xޘݛ�(���e���!n}y��Y�{'%s2�ew��@���'R�p��HM�e��Cҷ��e�ˇ�h��<�W�.�P�VZugG�Y�uS��ݏ1��𠛕!��L�ޙ�t��O�;>�z�*)=�*c>��3DdZ0o�vʓ��<��Ӭ.��\1F�5�ƍgR��r^��0� �8k>6s����]�!��	Ǹ�y85���~�h�Sü~���U��g��U-�e?�:�Z%�~kE#z��eU�e��������Ӟj��s �׊�8²u�8���=ON��t*�[P{C�#^v����V�/�בa��@IE�U���2�77�E��T���z��eU�e��������Ӟj�ܓj3:��ʨ�.��{2OoT���zV�p0�I#�r��8�EyF�8ơ�@IE�U����S8�����)�dMê�[��owђN�~��&�t�)�����n�p!!v*!��u���d���=A�2�S|���f?��� <ƍX�3�&-�=�&��誼V�d4Cm f�Lu�m�B�>�9��(�
t��Y�{'%s2�ew���5�"�r�7prEU�xm��"X��[���`m��O���U4��{2l���^���@�d�_C�VJ����̕���(��hG�U�Ƕ�2��c=�_R�N}�}����B�����8k>6s����]�!���)��ɖ�S7⸠z�V[�-jɸ����g����R.�C<�I��ZA���e6qR5L�/8'�G~+�3;��\���\��k�zph5)�� ��լ���MRs+-�rmE������ VU+I���_�����
; ��p*�����QK�>;?��Ϥk�;��|B}ø��y�w���H1��@�	��hN�q;�ǔ10\p c
N1�V&�����O�qTkή�Ádo�dvAg~�rk܀�#��˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F�;�sB*�1v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	��]���������ї4�z��pU6�M�S��2�{��΂Pkt����p���C��"�nT��z��uWU4y5=>F/ġ"���Չ-RW!�՗"$p\�>���S�w҄�^��(I�>'����	4T���\�nƨP�ʱ:��Ԩ�\�"ߗtl%�]Y�%���Ádo�d�x��u�5�h�br���lpda���?̕U�/j�g4A���{0Yafk��r.y����nL���~C�V�T��a׈Eg#f�z�q���<�{�!���"4��:@��o���KEd��]^X0��
x-	���'�$HgL��)������e��Q�Q&I`��=J'����r
���I}}3M�C,����|#^�Vn��l�M�c���=^��>D�c�lQ�����+�7끍J�[T�)��o�B��^�֌���<�a)�m�d�so�}a�C�ub;�;�濖n�P�������h=9.�Ύ8�qXF�����z�1�b$E�D_��G6il�٦p�d��r�b+ӄ�bİ��8 �����������c-�z��~��D:<^��`Y�F�����I��<�|��F+��4���LT K���Db�J��@��$L��%��Z��b,�A�zP��`�� ��D�F]�&��yJ��o�y��e����#"!��4DE'|�&�#�E�d��������y��Ld_&�Q���˛:���,�.ǯ3�4������$�A%q�
�$-���$73���'���))~�� ��-[�v:v�o���+����7X��U�?	r�����qˣ�ȭ�n�h�j�� ,� �M��U�RPkt����Ȩ�����orǟD�uiM���	�f�h�"أUMê�[��,�]��Κf=�Z~=���q}�w|�e��Fr	���Lz�U�pB�cm�ϒx��<��e��h���Z%2� r�BIWu�ׄЯxi��G\���L>��R��K)��x*�������ߘ�Ū�9؜�%�+���UA��́	P6�������&�E\׌N���ڪ���������&��᧲��\���L>��R��K)�|1������q�/y�u�?ƚ�z7���e)�A�?��R�%�vk��|Dm���v�@a��R���q�/�������x���hAklm�"&�Hb^�G���`L��U<��d[E�������iR����o�a`�"�X���-�+����S�_h�G�.]̌b;��時S�_h�G�.]̌ȷ�	����A+b��r�mR-AF\���L>�l�4��H��;.)iB��ve��Fr	�x�s]���uC#���3�`���U��A+b�펋��q�G�������?�?��(�G�l�4��H���ւ���z��Ă^�4�j�N�)�\x�s]���uC#����@�%/�w���j;&�PEMU�YGU���O�8c,}%@�s�a�`ھ�Y��^@!��?�y)����q�/~��:c�g���y�I�ވ௄㼤��sK�+�����C�������?�?��(�G�$�
�)���pL/���sK�+��q��j;w���ڪ����y��{W(l�4��H��?d��������>SELÕ�)X�J�$�R�n�KsFԙ�0e��Fr	�&�L4⭦�����.���"��	�x��<�����`B�)續\������kD2��)^>�b*b  �H�,3�V���C����?1�o��	d��p����ct��~wD[��8�Y��?��-7 �3�V���C�ۥ�	�VF-|��S��t��)�4������q�/L�U���;�A+b��`�,"�~&I^+������_����*�.ܓ/�(,��BpLÕ�)X�J�$�R�n�1���؄�
5���4�~wD[��@HK�OW�'n-i�& ܵz���K�ޛzṕ	P6���y��{W(l�4��H��g	Z��>�-7 �3�V���C��L��"܊VF-|��S��t��)f�]yD����q�/L�U���;�A+b���yy��z<I^+������_��������~,��BpLÕ�)X�J�$�R�n궓�rg���
5���4�~wD[���v ����W�'n-i�& ܵz�rApV�q5�́	P6���y��{W(l�4��H��bgz�Itt�-7 �3�V���C���?�VF-|��S��t��)���K��k����q�/L�U���;�A+b���g@+V�<!q�D�?�e�& ܵz��~��&����q�/N�߄�4�X�)Х��O@���`��n�[ �^�'���ߌ[R)Ms	[����Y`�^[�.(+��S�*���X��E�ސ�[�.(+��S�*���X�z�x��ol5v�I�D���t�:��m��
��\|��Ea+a�G3�u](⋼�1�n�,e����+8M��f��2R<�k{�����)�p*���n�,e�P���P����ӑ7�\�U j=�	"<�k{����Sc��6���y�=k^ŧM��ڪ�����4&ݞ9��h�xm��.�3���l��́	P6����4&ݞ9��h�xm��.�3���l�����q�/`�m0/���3�[U�Hl8�^L�a�E3t��,B���JS�gZ�瑪W¡����O�8HL�Ǳ��I� �c,�$��1�2>�1$�ۊb���`ܰ��ڪ����x�����jrk�PM娧�9�����B a�޶�oo=S�
J1!��]c��V�b�1�RR�,�*Ǚ62�,�X]t��m�.��H�c��1�U�)Qg���#��r�)6��9��xx�rDc��/�;��K�ߖ��klm�"&������r���aM"��r�F�*�_�JH�q���m�.��H�c��1�u�K|]���)ï�y0����;e5V�]C��%��Ob���q�/B%���O-�#���[��0c(��<>p����ct�q�p��k�_����m�.��H�c��1��;b��1�)S��#)J���l����+��2���ڪ����ݧG �ŴP��Cn**�8����>x��F�\.��0klm�"&������r���aM"��N�߄�4�X�)Х���qv�d��s���?�������r���aM"��L�U���;��n�^-.�T��s~���m!�X�����;e5V�]C��ؽMBW°��P'Q^|v���Q�cel��oW���V�b�1�RR�,�*Ǚ62�l�;�w���́	P6���ݧG �ŴP��Cn��g�K�
����QA\~���;A���g�R�"+�zN����!��ZB��M��7��@�7����A@h���X �Zj�����A�
��v�5��_ۑ;�0|������K�}i� f�Lu�mA�
��v�w�U�+8�yFZ�±��m>˟N�0D-~ж� ��%�B �n�6ӌ�Iۏ��*��Z�� �Q�c�,e(}� ��Z�!3^N��PMY(璪�cI��S}H�(���e��3�!`�mL��	���ـ�fH�k��j���V�2;��&������dMk�d�l�1�ԀUL�~�'Vb��1�pi�3h���X �{Ē�����B��+��р��U6�Q(Z����B�ip �-O���"h#�)��!��ZB��|��t�L�2�r�ēØ⭫�_(�!�/&�Jܰ�訑��3c/��!��DDxFp�}��GN�=�Da���BJܰ�訑��3c/��!�'�`�X}��GN�`��B�0w�Jܰ�訑��3c/��!lG�g�@rH��i�׻�L-�yC³n7^��_�۞h�G��+^zO��7�gI����I�}jn7^��_�۞h�G��8���7�gI����I�}jr0NA]��	�YI܁��(u���߈��7Y،��!��ZBc��5-?��_��cZ2TuFsY�w���*��Z����whk�_h���X � 6y�P�v����V�/h���X �=��[�U�EZj������B�>�9°e���)`� ��q&���1D����
�?<�!	b0�C}�,����۰d�����ca,E���d�����caQ��RU떐V�RDFR7��t��6�ǌ�lA�>P�2-i_e����͂���[ �����
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"pe�IC�_�\�����@J
A��w|�<��y�~/r�I��
����&�ɬ� VU+I��|�5y�n�ż2'�����ә�����/�4�}n'���a*�x���� ���t�ΊA�_i0{W�����\�.���yX�h���j�|�O�[���b�/���%H�$zȣc��- ��Ckӓ��_�d�dw.2�҇�L�Xڈ*-�kЄ�0v�7�m��=�c�}�"���}����{6���@�ȭ�n�h�9PV��'N\ǁٲ"q�Z˻r���5傟�����̝�wz�҄`�����'p�@�5傟������t_��?�e�[��G�^�,\ަ�It�� �Mx,�o�P2}�).;��L�O#t����n��]ߺ�`@t���@
�ђ�>S�8�d�����О.O��m�6$��\�v�ʁ�t+o����=ڏZ3C���BC?T�<o�nïi�q{�f��a�:&�>��s=wK��7�&d&(C�#�7#^�Vn�;ۂ��IÙ=�H7j�7'c���Hhqu!���5�Nn���4L"�+�va��2kYD���h�76AyW��t]g�LʛYoz?5��^_�V-��&'�ɀxmMê�[��s*)F����'n�^0o�J�%����U���"^ ��r<K����g~:�(���g��h���Ll�4��H���_�G��GJHn��z����̾���^�o�A�l>�0!Ed�yӘ�즤^9��-zS�YQ�l�h�76AyW��xTI��b�=<q>w	3��o=y�l_�F��)�1��bMI�����^ֻ����XP����.�/4w���BIWu��T!����
p��#�IÙ=�H�8��sb�����I�'�Tu��ek&}�tgX�a�Nڜ)�1��b��4z܂<��)^G�<�zL͊�q�����R�%6����8%Ǉ'�Tu��ek&}�tgX�a�Nڜ�D�&)%@��o� z��,~:��wJHn��z���hU��9�OZ+L�ʜ%�j@c���t�*�*�tsb��K�'�~ KB�~�.$(��A���/�������Qy����� {�y?k�[U���z-j>yR�_oN�h�����/�r`��\�vś��X&`�K��t���i�Oa�b��~��钏b�n���\���e�Q;���gq�IÙ=�HԹ��X��+ꕽ�F}Yi�n/�:y�0�6�]���~����_j���=���a����Wo��̗�����H��@Ő��t��[=U�Z硘�`�Jk�IT�f|��P�����ʜ耚ҵԼ�\�vŠ�B��닶O�t�&~f`D��>��5�i�8�
@TRsu�5�fT�9BDNq{�f��a�:&�>��s�N��b������y��Td^ I�2ŔE"Rbz ��ڡ�H��	��HY3���H5����Ęj2�B�[?T�K볋���B�|��t!�j8ZT'�_��z��̪��R�ë&�L4⭦	� hi��\�v�[�������Z���� G��`}��q5�ˉ�Įe��Fֻɬc��WNGMG�2�3�yc�A�̍~��lӟ����9/���`q.�YF�l�4��H���ւ���z�R[~�ҋ�zL͊�q��G�D�� �d�_C�VJ����̕9(�[�t1�e�BB�ݔ�]<̒�ދ"�@Ύ
+(ws��M�~�~.\ͦ�X��H�/gu`NT<��y��ON4�i-��,���-x×v�X�8����յ��\�v�]������_�sL�S|���f?��AJ��vNW�w��fD��o30�@C��iߗ�{�(s�O�+�t&p�10 @>$!�u�]aL�ɜ���F)��`��z � �o*�voj�N�)�\�[�!U��#:a�0$2�gD�����XP������<����Dg��y��tq�-[�v:v��I���w�����
�?<r��0��=�*��g�Ҙ�%Z_0@>$!�u�]aL�ɜ���F)��`��z � �o*�vo��sK�+�����C"���a����'n�^0o�+#�K>��{�TNJ?�s�E(��6�ג�Û��� �_C����3Yju�xߕV��n�N�������M�~�~.\ͦ�X��H�/gu`NT<��y��ON4�i-[04ͳ�����o�xɼ�\�v�]����:�ʟ�����R�fPذ�͹sC�MP������ܨ��+drV��,C%������&�I᳹L�@�2�M�I���ON4�i-y��{W(l�4��H��?d�����x�]�V���(c���^�����ܐ�!V��>�%�yZM�����k+�ZG��=�`#7l�;����C���1&&���O�耟օ�[[_rvNH��i�@^g��݀�����oQd�#��2Y���p.�����4���Zxgף�d��zL͊�q��G�D�� 㾨!zIDOⱶ��[U�˵�a��݌9�����
�ǫ�����^��J�Y�y��{W(l�4��H��q{�f��a�:&�>��sH�2Da���`�M7Э7l��A���ZL�4��L��Q<G�^���_%���}����Eڑi
�樄�ZWu)�=>�q�E#�U7�D�>���Y�J��W�y��{W(l�4��H���n@�b���U� ���_#8��shƻ9��[�>�q�E#�UJ�#��Iam�D6�U6qW�'n-i�& ܵz�?�o9P}71�9���9M/��:M/������;#���,�+V�RDFR7����_�b狡����
:�
5���4�~wD[��dk1�]��[GD@�F��q`E�cvR+G
WW�r>1�C�G��$���
G�|�!<��l�
Q:Õ�)X�J�$�R�n FA�׀��=���a�8q�O�4D��Y�Rsۅ�LT�(5�.>ؑ� q�.Pa�wI^+������_�����\��5�Dx�]�V�����TI��ԑ�g��@��C$����}��yoZ�P/�i;@��\q.�YF�L�U���;�A+b��@=��˓4 ؅��FJ��/��<Ӭ��k�K�ָ������Z�]�O�"�"m;��U��aVN�+�S��t��)���Owc�g��|����s�ݺᣄ��C�W#@-�ʳ87��Q7�j�!��>��&pR��a��\�}1�-7 �3�V���C���TZ�4];ˍH���@E�`�Aovj콙����x�w�.�/P���s ��5Ғ�>S�8�dy��{W(l�4��H���p�C����U� ���_#8��shƻ9��[�>�q�E#�UJ�#��Iam�D6�U6qW�'n-i�& ܵz��~��&�g��|����s�ݺᣄ��C�W#@-�ʳ87��Q7�j�!��>��&pR��a��\�}1�x���=�g,�5�TzS�@/{�&�q:i@_�8x<�A!ȵ��o�R��@�1�� G��ΜޜԽ/��O�[�.(+��S�*���Xw�߫�k�'���Xwd�n]Nٵ��_0��U}��s�'��U'j�0���XB�Uioέ���K�IE��q{�f��a�:&�>��s���V9̅����n�+�~�5:��f�~cG����`�o���PPV��ķ���4];ˍH��Oz��Z���;O��+�	6?�.�
oُ���O�	����'<�k{���� �g^M�va,�X����_�gD�����XP���-O/ [р$�c,�$��1�2>�1$��_w���<�UJHn��z��r9�3�<�/�1JpL�����ovr�8E�&g��|����rֈR�-�����
�#h��lNûL�x���hY�'�_��z�Ӎ�]��rň�����r���aM"��n�^���'n�^0o����SVc�m�.��H�c��1���ܫjc1��y���:M�b9���:&�>��s��]��rň�����r���aM"������GD@�F��q�b���V��]��rň�����r���aM"��^��J�Y�y��{W(3���P�٤\��X���XP���-O/ [р$B%���O-�#���[�"yd��N�}�g,�5�TzS�@/{�&q{�f��a�:&�>��s��]��rň�����r���aM"��L�U���;��n�^-.�T��s~�V�D���Kb���=���a��ږ�����V�b�1�RR�,�*Ǚ62�l�;�w���q{�f��a�sW��NZ�kj'�빔��D�.}���.D,����e!0�K�_3#ڸZ鎬�����r44���Y��sx��KK��~4"<��CA�}<8�� ��u��N�Y�N�rb<��z��}�0z�cUL���gM�6��㳧ٍg�p��HM�e��Cҷ��e�ˇ�h��<�W�.�P�.3�]���,J�l�/o"x�ȥR���z�G���h�b=m��2��o-�Qd�|��aK �!n}y��Y�{'%s2�ew���5�"�r�7prEU�xm��"X��[����fbK7͍��|��W&":��^�o�A��yoZ�P/o"x�ȥR���z�G\�}�-��q���K7�����8,�ņ�a�t���8���C���{l�f|��rs�i��=29��a)6��9��xx�rDc�ቩW<$��ߪ��wZ�n��[��{_8�Y��=�}�Vݨ7K������u��w1j��a]��R��$���^BT�ܘ�!ub�`,���1�@ �~)�sQ�I�0/zﴚƾ>�Cb�!n}y��p�VU��J}\�=�����^�o�A3��d,�K���C��jʭ��5���Ig`i�ҋX������S8�����)�d�R��K)����m+�q�g��U-�ee�@Rv����my$�N��lثl�;c��bW��7e��6ڿ �J�A����Oy���|���؀.����r����2uM�S�)37J*u�,�JL���Y�d�C��AJb�!��a]��R��f�Š,�8c<�@��_�igx��8�1�R@�e���ۧ} .�_���wg�!n}y��p�VU��J}\�=��Ӽ��2��}n	�Z^�t���,2����X�kX������`4�E%v�~������]�!���\B��V��PV�)ڶ�|ceJ�z��eU�e�����T�2���%,J�l�/]��-5L�S|��)����\�6�(�_3#ڸZ鎬����Ĺ#{�������犃�8�Qt�z��eU�e��������Dg��y��tqӴ����s��8�M���e���96��`��Лv�~������]�!���\B��Vjn.����Ϙ�J|�Qz��eU�e��������Dg��y��tqӴ����s��W�u��ó}����w�q��N���OG��_3#ڸZ鎬����Ĺ#{��2A���ϻ$�Zkԑ�]�Jg����-c �ЄW:l�mq���)�:;o�������=VU�����WΓ�Y�mݶ���č�Y���S�)37J*u�,�JL�������d)N�UE�B*�2���u���d���=A�2�S|���f?��� <���eW��H��ě�5/U�rQ��3c/��!`����J��<��z��}�<ͧ�:|C���m9�/s9}B�Ź��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,������[GL�����K+I�\�q��N��f�;�>)�~�`�0��|��].��'���Xw�����C��Z_�� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j����H��[n��B��X���WΓ�e'��ǩ����l�u+�v�~������]�!���\B��V�e9O��g��$y�z��eU�e��������Dg��y��tqӴ����s��~�̳o�"�D<�4_�;��	��Z\�i�æu�Q_�}{KS�)37J*u�,�JL�������d͇ :�s��]�Jg����-c �ЄW:l�mq���)�:;o�����p�ǔ|�b�ei�5/U�rQ��3c/��!w=����^<��z��}�<ͧ�:|C���m9�/�!������ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����&�2 ���������x��lV��(C6	�YI܁���!n}y��p�VU��J}\�=���T�<�����Z1~�g]�I���B��&���a�%�j@c�}������[
]&M��j���$5�}�����q>�~I� �_3#ڸZ鎬����Ĺ#{���Wl
% ��)ʒ�"��/8'�G~+�3;��\���\ ����@���d}�80�[X�b\g�8>!��J�0N�
���	�Bz���tU`f�g_3#ڸZ鎬�������(���R2�sW��t_-Z��T�\ �͘�f��p�b�z'hۉ)s���Ħ�q��Z1~�g]�I���B�龈4��G	������t4z��w���*#�IQ܋[���,d�܉-`�6�����Up��^��0� �8k>6s����]�!��	Ǹ�y85���~�h�Sü~���U��g��U-�e?�:�Z%�~kE#z��eU�e��������Ӟj��s �׊�8²u�8���=ON��t*�[P{C�#^r�3P���WT�j
�I��w��,�9���������a;�/8'�L
�2�Ot�ky����R� -�*3fN&����6��Ҡ��Nx]<	���rѮ�7]�8k>6s����]�!��	Ǹ�y85�ӓ��������@	Q��"X��[���`m��O���U4��{2l���^���@�d�_C�VJ����̕���(��hG�U�Ƕ�2��c=�_R�0��=��d�����caEyF�8ơ�@IE�U����S8�����)�dl�4��H���t_-Z��T�\ ��Sv[J�1ť�}<�&�/8'�G~+�3;��\���\��k�zph5)�� ��լ���MR�Ӝ�n����։�s/�yf��nͼ<�TD��x��3�]�����_�sL�jGC��w3�Z.��	.�V�~�-�r�e�L�]�തJ��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����Hg8l�6o���m�D��%�r �&M��y��Iۯ�oR���7�m��=�.U�m�M�L~΄gO�3f��*����f���,�LPkt�����q�s��D���e��o���1�^A���2y3���u�����!�|�{U���5����`K�8dn�����bū�R��_�}���\�v�Fp~�]���s�b�a��wq�,���Hb^�G��$~��������츕�)���~|K6�׍����}0�st&���\�v���T�©�����О.�8z����&��$�RmHX���׫�J��q{�f��aƨ:bN�t��n�ߒv0ܛ�	���8z���,�v���.�/'�����W;5B5Y+�Ȩ�� "��t���6��^hq��:@]�� �F�0��Ji%����hdZ0o�v��o!n�c����Q;�]��]!B���j�!n�x*4JHn��z��r9�3͌4s+�ny7ג�C-�;@���^ֻ����XP���E�z��6|ۂ��jǱlì��s��j�R�˼�\�v�?#<b��>
�5����`K��|I�"�, �z$���B�^ֻ����XP���3�Tt
�w|ۂ��jǱ��^J���F�!7��5q{�f��a��{oS���%�a�j��CK]� ������;ۂ��IÙ=�H��,z��Q;�]��]!B���j�Iſ�Κ+q{�f��aƥ��E\�����%�a�j��CK]���[�W��K���q{�f��a�h�T�����χU��3S���V���c�Fd�� �5����`K4���ϛփZ���0�JHn��z�~�+�oR��y�K3�(�C�b����M
3͌4s+�ny<۾���#?�o>��!`�u�!jJHn��z��nw=��K]��)H�bū�R잓��ǡX`h�-���K�vV��Mê�[���iz�2�Π�ur�͕`�Wr������	'���㳧ٍg��X����o����;e5V�]CSK�p��jO�����\���.�R���c&;ɋ��ă�s0�7��65�����{�#�^:��L-{����Nɋ��ă�s��y�TL6��W5�JA�;摼ڃN\ߤ��:���p*Y��Tq{�f��aƨ��T�f��)��}�OV��~�[_�"�o.(��"�K�b�Tn\���R���c&;2��6_�-N�V�R+������{�#�^:��L-{����N2��6_�-N�@�I����W5�JA�;摼ڃN\�#��ٔ��_�G��GJHn��z���[3fk���"q�ߺTZ94�&�v���D��lۍ���kR���c&;TJ�ov� ��03,���y�U�;fJHn��z��nw=��wJ?6�\�p!|T��c�w�V��R���c&;Z�瑪W¡����O�8HL�#OZS�5ǀ�#�^:��Le?�y�O��) �YR�3˭���߈�vJVt�l�褻�sv>P�^N2Z���%�a�����W-�PDRŔ�rUq��ɤa��)gΔc���г�IÙ=�Hd\�q[���B=>�6ѕ����;e5V�]C����gg˃�x�ZF���A+b����ʘ��"l�;�w����i����pRWl0E���n���7��5����`K�8H���b�"K$���~��j.o�c�\.U1+]�!�;$��|�ќ�T�0�q��I�&��������\|��Ea+a�G3�u]H�7��=B A�����>x��F�\�D�E�
ˮ��\�]\���e�Q�ԌN�����W5�JA���Q;�]�#Y;�9l?�u�Y�M�;e5V�]C���[���?S�*���X:�*��ܟ\I��:�;k����m~�?�x�&��{���l5v�I�D���t�:�(���\L�B%���O-�#���[�"yd��N�}�g,�5�TzS�@/{�&a7��:����%�a���q����g,�5�Tz�o b�ўw���Yl�B�rs�i�̚irZ%�� A�����>x��F�\��R�>�v,0=]^	�&Z�n��[���E����~��j.o���T�m�}�m7���e�;5�P����^���sL
�~�m��rp<�I�p\�WB����&�?&���2nv�J�IN�,\ަ�It�M:��2�,����|#^�Vn�^ֻ��!� c�"�;{
�js&,-RmHX���׫�J��q{�f��a��j9glg��`m��';��?2^�9<o�nïi�JHn��z�Pl��>YuI�H/�v��b�!cI�﹈�iq{�f��a�A����
�H�f���p.�������;��"-^ʆ�In��t,JQ���7γҬ�,;���ʘ��"l�;�w���;5B5Y+��A�DlO�
� �F�D0r➜~y��Y�I��;5B5Y+��A�DlO�{ƕ��w��\���\ ����@�!I/���P�>һo�%�ˏ8[$0��M"=� �n�ṘW�]��E�`�Աiux��#��V��W@0D�k�/8�-�'�����f`�g�W���?�y)�;5B5Y+� �i7�sp>�{ƕ��w��\���\ ����@�!I/���P�>һo�%�ˏ8[$0�����|w"�_%�C��~�&A��`�����i�t�<�<俇d(�D-rB}VGڝM����|%�[�!U��#:a�0$2RX+�/�o�IÙ=�H�&8���l�mq���)�:��j8HQ��e�z���V�RDFR7��ᚌ��J��:sS89�*uT?�Х |�8�}7E��O��O
+@~`��)�j�����x�d��v"n<�#Ƥ���y�I���re��BzL͊�q�� Ky��:~d�_C�VJ����̕9(�[�t1�e�BD&�t��х�NvV几���IL<����v@U?�_��B�e�D�*�Y�p�Yч���Ҟ�+����ɬ�@��> ����I�;ۂ��IÙ=�H�&8������5^�ł`?�孵����9�;�`)�,>��ve� ��w"iw4޴���`38��(�a�jj5+\�N<Wԭ	ƽ��~wD[����B<:��(�yudCi�[e���k�T��q��4�ͻs�	Õ�)X�JK�IE��q{�f��a��j9glg�H�2Da���`�M7Э7l��A���ZL�4��L��Q<G�^���_%���}����Eڑi
�樄�ZWu)�=>�q�E#�U7�D�>��`�H0����EW�փZ���0�jݭ�F���1�����h3;C$�-��qs�VY���ܴ�&�:�������͵���L�+�M�R��x���hA�q:i@_?�,�UP�`�P
5���'���ߌ[R)Ms	[��������4]���9r������Rm�Ƈ�hʨ}s����=Y��_�0z�cUL�����U��Qd�{�kGQ��l�4��H���^ֻ��!� c�"�;i^S$������7!W�F��F�<�:�9���P\S�Qo�${U��w�X�|0���KP�i�}F�sDE�:}|߿ v��>�uLC���+�$�-q�8��f��)d��y=�z��/
����X��Q\���-���4�5��?���q.�����'��Ӥ�nq�}F�sDE�:�]ƭ��&��}g��u"��*�ΊJ~��ڹ 	��\�v�,JQ�����3"��0�;e5V�]C��( _��}mAb�+!� c�"�;���j��1�RR�,�*Ǚ62嫗���}�8��f��)�b���Vx���1�|�c��1��;b��1�)S��#)J���l���\�M�u#RRJHn��z��r9�3|�bІ��xx�rDc�5��ja~��j.o�c�\.U1+]�!�;$��|��XP���i^S$��1�RR�,�*Ǚ62�y��{W(3���P�5��$�/vD���?a�s�ݺᣄ��D`�%�����r���aM"�������4��5���R3�A�DlO���=��s*c�r�w����bU^�u���d��CE�-�EU��P�:^�J�_-�_3#ڸZ鎬����b���h�6jK�:[f��,2�����^���@�M�{Z$~ҝ~�k���M��������}����� ����+������!n}y���q���U��ED0 � ���ѡ�e�LZ\^��[R�5z���t�|��].��'���Xw0X�����!'lBv}���S9w�|�&oA�\ֆa��M(��*��w
j$�(/�W���?ᵏ�q(�܄��� M�č�Y���S�)37J*u'H?�׳�#\�)�`"8M�.�<���!n}y���q���U��֎)A=�s��]b_3#ڸZ鎬����8�������F�!���Fi����o_3#ڸZ鎬����r�1�	�0<�x����am��%��{l�f|�ό���.�41�(�6c�s��]b_3#ڸZ鎬������yA�'F�e!0�K�_3#ڸZ鎬������Wr��a��9/���`���6jI�־�2�h�ˏ8[$0���V�2K2S�)37J*uc�A�L'M�Kc�Iؿ@I�I���1O�~oua(􆿳�ʨ�6�j��2+i�27�yӘ�즤��`3���j�w M��b�M%:p^�vi|���؀.ņ�a�t���p
��9�-M����S�)37J*u�v3���?���XM���ӮY�E�63X����8!�T�vdWS�讒 �����'^C~o��Je�Bmy;;���0��0��}�<l^���f�]�!��	Ǹ�y85��NÍ@�xx�rDc�O��Юlb�Ȯ��ߊ�Г�������zl)BO�>	���n�sӠ�k-q�o"x�ȥ����\���ݨ(��y]5t��v_3#ڸZ鎬�����r44�����6�z�
^������E�]�qw?����
�?<�N*��;_3#ڸZ鎬����fS�gG8��7��~�)�p�=A։�Xs ������>q'i<c�!�΄,�H'u$��U��{\>����Y�cӴ�"�6j���'��mr<�ҋX����0�a1i~JK>��{�T��p;��$�F#I�%�[���69[̰�&��YcH���V�B�_�+�)��� Y�b�7��S�:I��w��,����8d��'�E�Jg�S�(��ɒ���9�dMbZ鎬����C��5t(�/���jbPhrK�@<,у7G#+��Q2�+�Y�-�H[����>�h$G����%y���TD��ό���.�"���0Yp <�r�\�EyF�8ơ�@IE�U����S8���Z�/������i��BT�^��a(􆿳�����|�z� �߳G!�a�`��}��(�
t��Y�{'%s=ͱu���b�% ���X��������`y������3'�L��ߺ2���;=z�z7G#+�Ǘ0z�cUL���� @c�8���/�3�;��x�� h�",oMG~�/��;`5/�I��w��,c�A�L'V帧���W¡����O�8HL�*��T�����`y�����u��Ѷ[?4���R;W&�]�ר�TD���9�,�w�8qTmI(xe�0
A����� �|x���� ��X����(h�š�b)-�uA^�Koْl��]�Bo�;�>8B�I:׷�F����������Ψ��F�x`��:�,�qo�,ܛ�	���J��p;�a9��Ў�4�t=�j�.�/'��Y�
Q���n�\�
k�#2��I=�=�l�Lɼ�Q���n�\��	��u��t^ꦤ0�7��65�\�c)rJS](������u�|z�$��e�X�+� �{�c�vI��?�-� ����w)��O;3<�U�C��z����7��j�5��iagƪ��U� ���_�L�;��G�GK�\�Ԁ0}�����Z鎬�����ꢃ9@;�1f8i,�#S�)37J*u)T{6T'�9��8�'�Z鎬������v�R����kK&�h�]Z鎬��������e)FC���� ��_Lj7�4Z鎬����SkRH?)ř�b܉���8��a�R�S�)37J*u)T{6T'-8W,UV�TD���rs�i�� ��*b��g���ޔ�owђN�~R�wX��j�jz+ ^���j��fj�TD��ό���.�Dk��v�Av�X��s$��2����S�)37J*uc�A�L'�H�N�P]��Z���Ga(􆿳�e�&���6/����p����N���5'���Xw�j�7��o�${U��w�X�|0���ߪ��w�������8]��?L��we�ÄҋX����@�ڗe'�ح(��A��	�_�*�'�D��q���U��G=X����"�f8dP�!�c�餯���Z鎬�������(����T�3,��BT�^��o�${U��w�X�|0��X��������`y���13�3��ŧ���X� E���K6,I��w��,c�A�L'�}�4?k�a��0�BE�9Y}��P�^�V]��}R�wX��)s[�3��k������餯���Z鎬�������(����������TZ94��h���o�8���/�*l�\:6�
�\�W�EC�2[QvA�m��w���Z鎬�������(����������TZ94��h���o�8���/�g�y�ޥ-ju�u[�z��-���a@IE�U��@�ڗe'<y�׀%\��߸^`��TD��ό���.��N}�}����1�G�Qc�k]m���6�vg;Je'���Xw�j�7��`�|��K�z�Wǖg3ȓ8���/�*l�\:6�
J���o3c�-��;�����!�!7��TD���rs�i�� ��*b��g���ޔ�owђN�~R�wX��ɞJ$��^�5M�YYroE�4rh��|� ���]�!��Zˎ�f+[O��ɔ�<5���3�n��#��@IE�U��z�г4>\��p}�	��D܂�A�ϑ��[��0Q���g�ƙi�Hύ|xy��"����S�;Fuu�p�w4�i�5�d��-��?�z7����b���1�߽K}��׍����}0�st&���\�vūx`��:�,�qo�,ܛ�	��|��	(���zL͊�q���19TH��@���U@���:��F���V!���IÙ=�H�^,|���Q��t:(� �>u;YW���\�v�ȃ��X����+���e����ȇ_���ˎ)&�E\�w`�|��K�z��5��8�t��\�vŭ���z��2U\���\8�ǔ4�_a�CK�H���Վ�(���k�N�� �\	��rR��^ֻ���(_�<���Iۣ<�;�'��-d�Ry��\�v�w5��\�p!|T��W�F��F�N��B�)Y�	s��N���:�?�_�G��GJHn��z�dD�J'/��ڧZ��7����.C�M��LG��j_ R��L���+��g�ڧZ��7��M�P�Wݣ�Tǉl#�'�U(�M�z��IL���M�U2��IY`���@�~r6(�睽_���wg�|��].��'���XwM��.��^."�^�ѥ�"���$v�~������]�!�����#e;7mg�oc�.[K��m��/��*�, h�r_3#ڸZ鎬����b���h�6ϸ�Q�E�DMP˞+��Y���?��;�x����������Pma���n��)\���M�^4/��?Ev�~������]�!��3P1������c�v�ߖs��]b�|��].��'���Xw�$
�Z[��ck�Bɉ���o_3#ڸZ鎬�������#�2�F��M@3%�w����$ĄҋX����@�ڗe'�0]���!Vf����aU�7L�<��z��}�Q2�+�Y�W�!�
���L��Z�N3�L�t��n�|��].��'���Xwd�n]N�}/A;T�c�owђN�~��&�t�)���y��lDY3!�buh�A �sbZ1~�g]�b��T�Q5��P�J�W��Ws��>�C�~�rѮ�7]��!n}y��Y�{'%s2�ew��fpx��p��HM�e��`y����G=X���Y�����Y'b�'=�(_��Ym�@%7G#+�Ǘ0z�cUL�JJ�4(o�a\Y�����BT�^��a(􆿳�e�&���6��&���'b�'=�(_��Ym�@%7G#+�Ǘ0z�cUL��W?vxb�k�N�� �\	��rR�^�V]��}R�wX��W��+�}�5D��0h\Ef�>yf��i��]�!��.��H�=�N}�}����1�G�Qc�k]m���|��].��'���Xw�j�7���|��{�r�\	��rR�^�V]��}R�wX��a�;�f����X��֑xGV���	��� �S�)37J*uc�A�L'�t�N)�~T-��qs�VY���/7R�%�T�\ �͛A�M����0Q���g
3K������rg�D7�ҋX�����=�슶}.�Q�º�F����U��~T������+GkۯΔ��Ig��ĕ;Ø݅ VU+I��(�@$.>��K����\#+��Sз��x��@���U@���:��F�ʳ�A~�0 �i7�sp>4��D��6`V-u9�`�q{�f��a�J��Ԋc���R��K)�n6�"�j�-�l���n�2��`���\��G��
�OU:�d}�n4$����P���{ƨ�X�*�7>����p�*_�v�~������]�!��	Ǹ�y85����Z�m ��ߪ��w������Y�mYj'v�~������]�!��,��灋O�N?c�<��6�|��].��'���Xw�9�RL6���nf|FN�!n}y���q���U�Bă�CL��Ig`i�ҋX����@�ڗe'K@4I_�GZ_3#ڸZ鎬�����T��`S�������{l�f|�ό���.��5XsGf�בa��@IE�U��w�B[��lQ�$�k\_x���� �~��Z2��rtK13��\� VU+I��ƴ��������W��x�����+�@{fT�1�߽K}��׍����}0�st&���\�vūx`��:�,�qo�,ܛ�	��|��	(���zL͊�q���19TH��@���U@���:��F���V!���IÙ=�H�C&�����}�K�
�4l�(���.YT;�u.Z鎬�����D�Kw��L�?��
�Z鎬������p���ȥ��9�dMbZ鎬�����W-O4�؏�F����U��~T����Q�41�&�0x ��lzb֡�ɰ�s�!^�l��^E��fi���K�Q�����R]Y�~�����Z鎬����D���Ru�C��I�"j9�c�;J���C�<�f�|ߐ=�%��)�@���e�cNơ�&Y��V�c�	��}����ܴ/a[B�����'���Xw�p\�p���"2�#�>��~���1��B����qC�<��1���?�{�W~�_3�mE�_s���R�AZ鎬��������}������$h��qa]�݊3�D�A[�rd�׎o�|MԲ����ﻋ-���C�M��N�ۥ��N��>�S�,֍�Sx�lޞ�ό���.��
�-�������ɨ�ML�9࡯�d�٣�����6>���]�B��[S�7P��T��]�!���1����m���!�����Ig`iZ鎬����Y�V��#qa��w��[B�����'���Xwa'�<� \��x��+jMf���9���q���U�pzl��a��\�(Ƭ;1Mf���9���q���U�f��'����Oy��������
��#���	�U��*}��L����� �P�b���l�;�w���=e��i�W+`�x�o���{����4�u>�[�9q�Y�{'%s2�ew��� �GQ鍚p��%�g��U-�e5��e6²*�wX8���R�Xe����>S��J�"�T<L��P�b���l�;�w�����?�����qi�á[�6���l �����4���ʽ�n8`ݧG �Ŵ
"4F��l���D��q&��k�S��g��U-�eoC]�<9�v'�P*�cz1�� ����Jm�W%�s�I�5�,���'�f#�}N9�h�Hx�D,�d;vt����3Y���6�I�{�IQ{�50�Vr�N��+�4�֧��L�q����Q~��:��'���Xw�j�7���F�xE�W`�|��K�z�Wǖg3ȓ8���/�a'�<� \%5�Ψ-��;����Pn<��Y(�v�]�!��	Ǹ�y85���t����?�o>�:�
���O�g��U-�e5��e6²�KU�����1�G�Qc,e(}���=Y��_Q2�+�Y��)�`E5�'�r��'q2I������y����*0oό���.���K�Q�Y�����Y'b�'=�(_��Ym�@%Z鎬�������(�����"��a\Y����t_-Z��T�\ ���|.�Tӏˢ���[�� œ�Ęlz������ﻋ-�����S8��$�DB��H�e�X�+� �{�c�vI�ߪ��w�������)�`E5��{�^�X�5D��0h��P
Z鎬�������(����mA�������b�x��+�p�U�C��z��
������y��ٓA��ɜ�\��R�wX����K�Q��&���q�GR�W&�]�ר�]�!��	Ǹ�y85�i /�?���ڧZ��7�ߪ��w������$Y��C�
! R�7��1�G�Qc�k]m���ﻋ-�����S8��$�DB��H�|��{�r�\	��rR���"X��[�z�C������ıψ�I*�?��m�±��m|�qF)�('���Xw�j�7���F�xE�W`�|��K�z�Wǖg3ȓ8���/�a'�<� \�����$#ZƧe7��
`����0�E>��=Y��_Q2�+�Y��)�`E5��{�^�X�R.p���M�aQ�q���U�pzl��a��&5�/h�� �����k�~��Z鎬����D^Rm�	�0i���WX|M���k��s�KT�n~�x�����&�EȘ87Yxe�ﻋ-�����S8�����)�d{[���G����"X��[�{Ro�č�h߹5�(��N�g�dez��w����yoZ�P/2�cQ皃3�I�5:��.@���K�Q����
�?<J�!�Ӑ�JR����]�!�������͋{�p㘂��5��4`U�j�d�|�T�bj�V�c�f�:3b���qq���"�Ee�6;�ﻋ-����2�77�E9g�M�G�n��| �u����@ ��S�0/������;��\�?D�>*���!����|w:J�d�٣���9�����!��I\+�8@ͻh�C�E� ���s.��n}7���qOΛ���[=�@��r�UHK��q���U�]���V��+$OF>�X�}��z�?����ra��pzl��a��>�u��8!��=e����$J�LPkF{������%Hlܰ�|�)n����S��m�1T��jF3�$��3�M��.!y3�Jp����a{ΨmZ�az�6TrDE�#d��!�d�٣��c�A�L'�f?S�$�R�n,�	�X��;"��PÛ��+�p��
��gl�4��H�������4��Q9�5��5��`y���pzl��a��B�M�5����a�|��52��n2�d�٣���9�����LL�ΌqYF��J���"��#��b�N3��E��RQn�';�=��6�p��xi�[�=�5x�=�r��R�.����]�!��b�#lx0�߫�-H�/�L�)�y��Z`���U�ZG��}ݓ��E�i�T����n�Y?v�<�d�٣��V��4���;w>`�2�o�M�{���'C`ø����na�Eb뾯��g`����^E��fi���K�Q�b��o�I�z��a7��ﻋ-����2�77�E۾S���*�[�·��`נ�%���L;S���s�����k��&�8Z鎬�������(���osl$й���&���WX��y�g��U-�e?�:�Z%wƄ�{Ƨ\�$�������\=����2w�7H$�DZ� �T�٥��T8j�Y��!P���b6H�W�^}�-y�[�P��n��7�Sx�lޞ�ό���.���K�Qs@�&eVC�8M�.�<��ﻋ-���C�M��N���H2�)�؁�u��m,3���-�$��]�!���1����m/�n�*���$wc|�fw����$�Z鎬����Y�V��#q\k�{j�$�u��m,3���-�$��]�!���1����m�ρ;C��f������s��]b��=Y��_Q2�+�Y�ݓ��E��xsթ��� ��M�d�٣�����6>��b02�O�x����am��%�d�٣�����6>��T����{�M���5^sȘ87Yxe�ﻋ-�����S8��y��Ʈ*M�����^�V]��}R�wX��8����oo��u&��P�:}ϼ 8�������*�E��M@3%�����B�['���Xw��t6Qƹ)5�(���{�eV��0�dy��8ۦ� ~�p��XөF�?�y��h>7�*~}�_n��իe�4�r��n�"���:��-�3�T�Ҹ�X�y��m�Y��E�&����f��jv�!d*�[���m}����X�>P�2-i_�d�Wz|��$��4[�l�zq�����Z���%;_{�& �^�͘��r��T�s�6�Hh�4l6���Fc���LV��f!�A&�c����)t&���J`���f��0���E0)�BoE0'�fg탷�J1g�J�6�̺&?�N0)�BoE0'�fg탷�J1g�J�"��?^0)�BoE0'�fg��mQL��x��M���N��0)�BoE0'�fg�m��3xȀ��aI�V}P0)�BoE0'�fg�m��3xȀ���M �})�}�����T��.��W����u\��W�7"�I_$\�j�V��v�@�M�¸mA<�SNp>��Fc���L#*ު�^��J�Y��.�u���M^!�3%J�/�x�/7H$�DZ� pzl��a�S"#T�Q2%M��Sx�lޞ�ό���.���K�Q�h�6Q�7�0ʓY+��Sx�lޞ�ό���.���K�Q	W��^$k�i�kL�5N�ﻋ-���C�M��N��)v��Uk\���eq(1p <�r�\��Q3U�eT(�q���U�pzl��a�S���^RSŞ�Ӣ�Mf���9��Y�{'%s=ͱu���ɋ��ă�s0�7��65��Wǖg3ȓ8���/�a'�<� \[�	m�KԠ��ͩ^��Sx�lޞ��rs�i�̚irZ%��<�k{�����Wǖg3ȓ8���/�a'�<� \[�	m�K�3W�ǡ¶֢��s�K�� f[�rU�Y�{'%s=ͱu���ɋ��ă�s0�7��65��Wǖg3ȓ8���/��Î+,�C��XK�ӻl���r��V�6IWJE�a�1�H!�O��['����owђN�~vT�V��|�������c�A�L'�f?So�${U��w�X�|0���ߪ��w������ݓ��E�� �߳G!vA9�,V>d?
�����="��x8I���l2B:���XK�ӻlG~1��v��pzl��a����L�Y&U%����f�Mf���9��Y�{'%s=ͱu���2��6_�-N�V�R+���Wǖg3ȓ8���/�a'�<� \[�	m�K�P�!�c�!�}�"Am�.J)���rs�i�̚irZ%��ߤ��:��*�I��p��HM�e��`y���pzl��a����L�Y&�yO�6iSx�lޞ��rs�i�̚irZ%��/�rŗ���zl���yp��HM�e��`y���pzl��a����L�Y&E�̜��W�1��?\��ﻋ-�����S8��$�DB��Ho�${U��w�X�|0���ߪ��w������$Y��C�(����D��Z��_��Ym�@%Z鎬�������(����o�F�\���e�Q�mƿ�Lg�g��U-�e5��e6²�!`���� f�Lu�m�k]m����5�ź�ﻋ-�����S8��$�DB��Ho�${U��w�X�|0���ߪ��w������5�e`��9�<X��u���zW�'0+��=Y��_Q2�+�Y�5�e`��9�<X��u� �>;V���_���ݢ��d�٣�����6>��zK��i�� ����*��<[�+ꔏZ鎬����Y�V��#q��p��m��0Y d��M'�F2����=Y��_Q2�+�Y�kѶ���� �}r�HDʞ�sB�_�	�/��]�!���1����mφU��óv~�z�xE�?F ����Sx�lޞ�ό���.���K�Q����/�4n�Y?v�<�d�٣��c�A�L'؄�f�?�&3�-��_�owђN�~R�wX����K�Q����
�?<.���6���(O,[ǘq���U�pzl��a�9g�M�G�nE�̜��W����u�u��=Y��_�0z�cUL���a����"q�ߺTZ94��owђN�~R�wX����K�Q�	y��J��U%����f�E�̜��W����u�u��=Y��_�0z�cUL���a����"q�ߺTZ94��owђN�~R�wX����K�Q��Q8� Lڈ�|�Mf���9���q���U�pzl��a��yu>I���mϘ�=Y��_�0z�cUL���a���c,�$��1�2>�1$��s���S��*��Tɀ�X���A�L�m�M�����@�i;2��6_�-N�V�R+���Wǖg3ȓ8���/�a'�<� \�]VI��Z������D����R�AZ鎬����Y�V��#qˢ���[�����&�D4�ky��ﻋ-���C�M��N��+w�7�P�a�⏡�uܲ�?�t��d�٣�����6>��-r�^�Q�<��A���Mf���9��Y�{'%s�
>���j|~��A:�
���O�g��U-�e�t���R���ıψd�����ca����{�/��=Y��_Q2�+�Y��׎o�|��։�s/�H�c�D��z��"?#f'���Xw�����U�/	��Ɛ�dN+xޔ$c�����FK��)�H����[[��
fD����B�8r\V����p^����.����Z鎬����Ĺ#{��a'�<� \�/刲�Z��F<-č��_��'���Xwa'�<� \���B�F�[B�����'���Xwa'�<� \�\7���#I6�q�3)a�d�V�Z鎬����Y�V��#qz(�j��Td��p'k��o��`��[J�	���3�rs�i�̚irZ%�ސ�NJ/��!�#��W+Δ}M��R���V�'���:y�g��U-�e5��e6²"x��@׋8FZ�±��m0�t���M/	�~�Z鎬�����"I�����sy�������D��ܒ2W��4�`#������^�
�CӞDvp<����[�O���XS=��=Y��_�0z�cUL���a��Mê�[����@�nf�����r���aM"��r�F�*�_�ņ]�yk���`y���pzl��a�7�u��\<�m����H"Sx�lޞ�ό���.���K�QM��EכPT922�d�b҄cA�]�!���:�o��d���d�o�P2}�).;��L�O#t����n��y,d��6{a�t P�^�\MGl�<���{��ZT��6|�� =��_�Z�G�a}Cfx��V$�w�Wή�li|��Q"}Hi���#2�}����[��Y-��J��׍���
�6���.�H��7TB�7a	�����Y�
��3��X1�'�3�$ �#^�Vn@j�cq9��M��0�d�Sd��_�a���n�|W#"���vL�
; ���<����z��ɧ���7�)a���%}D������h�br���lpda���\��6m��B��${��?�J�Z��]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gV��Vv;�Oe�d�#���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂Pkt����p���C����s�x�9��喐Hj�Y�_�]	5r��ǃ����_����~#�\��OA�z޷S�xo Y�B��
�M�n����x5=��{t_�sVh�a�|�&�#�E�d���������|��=;��|B����?�IX[��O2 7�,�)�C�BS��g\��ı�ZnZ���qq�c�@,��ڬ�A ������ĎɌ�[9�-�Ҧ�{b�J��@��$L��%��Z��b,�0g���>a��v�<�RohWt�_a�fC��0��:Y����i%��ό�;�LȫԷ�/��Ϥk�;��|B}ø��y�w8#�RC�G�G~��6d��R-��2�����Vc2�����VcREBR�hHr�A��5�V�����w)К��g: k��2�����Vc2�����Vc�vA�1lX�c�M��;�3���v(p$�/B��t��!�,*}q��@��7� �B<=OU�۞h�G�G��} 5s��;�H���o�#2�	n�����0����T�'��x���ͩ�Z�K��{q�E�ـL��u�d�!�{�x�173��i��.;߱�-(��}b�ꎜ��t���]bC�I�š�h7�a��c�,�[`���!i��J��y��ݼƐ:�`���I�&�``��B�0w��[��U�D���L�b3NM�d��_��;�H���o��l�u+��[��U�D���L�b3NC�9mE_ݧ�f�;�>)�M�?��?+�r��`����s7b`?�'n��c�,�[`�t���iqFEĈ�d�1r6y_s� ��DZܤ�jh"r��c,W� K91j�L�uVB1��0�캧xӍ.��L-�yC³c,W� K91j�L�uVB+�o'���<���I�&�`E�b�.�.oA!�?2���-�)d�7v?�[��\n��*^������O��K�\|��Ea+a�G3�u]˴�����x_��s�֙���2A �����qOΛ���[=�@�8�'��Tn��Ո�Q�6�yP��C��?�zٰ��A6j�"Hs"� ���k�[�Ɍ㕉p4���\�j��fxB �y��	��e��Żl5v�I�D���t�:��Zcqe�+�;��|B��}zϹ#�H����.^݂�`� t�*hH����.^T�3w�?�D����\�V��	��yo��Rn��$7E����QS9�<�d���Q�^�� H$[4D���Ӻ��L�~�y�ю�?������I�����5�2D�3����h��=@ۜM��0�d(_\�^?'qKy���\N}zp�jN���xX0A.��(t�	��i|Stߛc�-�}��a��E�ȴ�T)�9\�V���$73���'���)��"�$��7��s�a�`ھ�D0r➜~y�wR�� �K�C����t�8���l�4��H���ւ���z�ktr[�h���̋8��s�$�R�n�m.�>"���(K�&)�*C�8؉b�'��(�~��e�.5�����O੺���N6�A{d�F���,c0�2�������>���F���<�B6Ji����A{d�F����`���u�r�S�<h'�4�!R$/���d}��[�ƭM^K�?�."�7���� o��e�D�$�gꈺ�x\e�L���8T	��sK���3M�55^��7���^Bm�m���Ыl���aWg�D���Sl�J��G��Ӽ�ʞC�ݢ�Iv
����Lc�TH������7���I�L�D�u!뼤Ÿg8V#��4�x&ʕ#;���{^���B%���O-�#���[�t
ZZK�z�f����ֹըQ��kGQ��l�4��H��x�d��cɁ#g�k��`�
}:�������]��:s+���j\�ʤ�/�V��	��y�@�3-dns`&Ѡ _;��i�1Sx�F?���-�z���ԿK�^���c�i	��e��Ż)6��9��xx�rDcѴ��B�66��ѵ���mm�Ҟ~N�����5�2D�3����h{d � J{?�d���&���h�p3B���X0�ޛ_�.��%��v�ځc����]ԟ~�[-���X0�6�4q̆8:F�c4�JE�{�F�S�ǧs6�6�+"�{!|�+�������gh���u�![1������R�E�M�b!yM�ڿ^�$��o���Ja6��>Y�B�5�]�i�r��y{�הr�=O������M@3%�e)6�_X��E�+kg(S��^7=k�Rm���0��� F*,ƌN�jK�I�q������/f.������H/Q����I�3" E���M@3%�9tJ/.�HL���dL7A�k�6�жD�n����Wa-�>�ТKH�{?�7��|�Ks���Y�"GF"��) �lQV�Z2�M�Q��y]�/HT�Y�[V��M*�x��<�����`B�)續\����'ò�������?��Q�&{��8�a�;"��PÛ˻Q�0+�k���R�bv=��`x�¶J1�j�A�i�A��Wa-�>�ТKH�{?�Us��'
��T���x�;	㯰�׏�����M��ܐ�}�ё����x���X�����xp�"�/�B�M�5��Z}��_��
wc�l�4��H���F(�E���;�
%�����DRŔ�rUq��ɤa��)gΔc�>�#��FY���$ �'ب�ϗ&P ,��rQ��s�����W��Qo�X3,���h��ۜ�����S���o�F�\���e�Q��8zK��	N�h���
�m��ט��+�p�U�C��z����7��j�5 )��\���,�	���pg^���\�}���d���Z�B�dhf"�������d���X�����K[ҩ:�y��$�R�n,�	�X��;"��PÛ��+�p��
��gl�4��H�������4���Q�V#��� X����Y^8�����D����^V��	��y=Aa�PZd}���d�l÷{H�D�p��M��HSq	��8�z�-��o�${U��w�$Q^ǐF����[u@�59����ֹըQ�ݧG �ŴP��CnxPT����L��S7-�;��|B݄�$`�ڹ�"�j�f��gFĝ��̡L��)�Iv=��`x�¶J1�j��5�"�r�~G��;ؔ��r�C���$�&V�B%���O|�3�d(]�/{��l�ƶ�~b�!j���.Լ�;��|B��q*(*�6�i�l`@��Z,r�_�n��j�=4ϋ[Rc�I;b�6mb!��u�t��D0���0�N�6e4����e�0
A���C���s��A��ˮ���o�u�/�ge��u$ħ��(vP�T���ol����/�?|�z�͉"_� N��r*$7�门Q��Ȝx�3�ס��wH/Q�����܄��� M��v/�ED�O��Gy7A�k�6���6k���$��M�W8߸��S�Ȍ��O�D	�%vF/�-B	y��3vQ!�3��hi�i�����a�s+���!���2o$�]��9�GKP�2�����Vc2�����Vcl��w&� 	���#�|"ap�� s;���*5���(ZH4~��2�����Vc2�����Vc.�
͹U�X�q�	���t7�j�.�q&Ѱ��Z����e�D�"fwJ�yf퀔������	-$ߔ���e�cN��M�� Qp���u%#��vWT�{�Jv�~g��?L�63@(4Pc��?@W���lC������J%��ό�;�LȫԷ�/6�����n�{5�G�<FJ�����Z��M�������"X��[�^ǣ�,Q�!�'��C�#�˛m#%��짐�CY
-����hB?�F�n���V���Z�4b����*]�?D�>*�o�g�`G��Ϲ-����M@3%�� o���YdZ0o�v��?B����ߍ���������ri���w9���I A6˃rG_�f����4��yq����ҙ�a	�lì��s�w.���%\�)�`"C�#�˛m#%��짐�CY
-����hB?�F�n��>7n���`��Fi
uS�4q�
; ��#f(Y��[�n�{5�aX��;�x��B#ݧ{0�(�G#��ӆL5��J; ��#f(Y��[�n�{5�aX��;�x��G2<��\�t]�sj�yIZC�#�˛m#%��짐�CY
-����hB?�F�����Qw'/֭FӸt���(�x�@�
�����;��K�"Pc��?@W� �!�3���|I�"�,b��:ՔX�.�	�5���#�^h-�(����C�#�˛m#�9��^K��9�)h�A�pS9�<�d��p�v�J�W�g���0������q9+t�}�T*@�F+��x��H��}c	��e��Żl5v�I�D���t�:��s8b�.��;��|B��W��$~�D�;E����� p��3ZW`����7A�k�6��9R�$P|g��D��l��z�͉"_�����������Cᣨ* �|O�ܩR����󀼍�M��7�&�(���D,���s�Mzr���Ƣ)ʫ��6o�]%����n~�/=�}{&�2ĥ)���� q�.Pa�w�8��M9B����*�E��M@3%��H��	W� OLfq�n���&�E�΀��h���,��5�Q,�=��1aԽX�t����g!4�s�8狗嫎�r��<Н�H��	W�p4�Q��������$s7A�k�6��I�ߋ��خ�&`ӌnA���qa���qOΛ�ٰG`ey,����N=��ΥT�tJ�1����ݾ-/�uu��ڿ$�)�vxe�zA��;��|B]it7O� �a�� �ό���.�j.�0w�q�g�
"^߫��.b:��8�z�-���kGQ��l�4��H���0�0�h��#g�k���g�0�u!��I\+��o���9B<0������q9+t�}@[�_zβrꢯ�wv�� ��g���]~�7i�@h�3�k�2�����Vc2�����Vc2�����Vc:'��β�=7B����ݟ�9��zԔ��_�c�Kʻ(ZH4~��2�����Vc2�����Vc2�����Vc�6=b�m.C6w���8��ͤ	j�e8�m��ِ�o30�@C7��G���ږ�3xZV����k,i�OL�JP�1z�:맷&�������P{��^��B�t�T�/7H~s��S=1�0������Q�h`9�ӳ.�c�'�\F��.�>�?��~g��$h�`+���7�ݒ}dZ0o�vʻ�3]r}�/�/_��qĞ�#�1RdG�y#�
z���)x?3ᇔ͔Ci+v_����k� ɮ�iW�X{����?��~g�5t�&��f�&�H�`b�h��8Њ�&g�ŏF��b�^jEml �t��61&E�۾t�V�t�:�c��1���p�H	�v�F#�5��*3M�АY�Q%~��2xJg2���fZC�:Gv��^
6��g�dO�9��9��7��7��W`���~�^H��DX�2�o��ZU.6�-�T��i~U�������A���/GU��3�y[�g$\�]�77:�2࿦7>�-��F�YM%����.�b��ѳ��|ai�>�
���w%f�������l+�%��v_���W˝�ѷG*p�[�B0�iY�<*��âcWx����e�(��F��� �8 �\ aNI�iǆ5%�5d���y���W�y�kv> ���ٲ/1NF���ݰu���3K�<�H%�'a��b|�No�{�׆lwhl�F�[��)��孱�������z�{� ْl��]�Bc�jv�Тk1�%n�@��V�����<o�nïi��PL{�ϰ>D�c�lQ�(��Q|3��'�3�$ �#^�Vn�����'MRmHX���y�XZ@po�ͫ��;���^hq��:�V��ÑR ����*��Y~��`�J�(��Q|3��$�R�n�9j�ʛ�́	P6���$�R�n�6Knr�7γҬ�,;Ot�@G�,�29a���Q�[<��Md���Lz�U�p��(��ʓ$�R�n�m.�>"��F��*O��5�"�r�x×v�X���0�F*�ZM����|%x�s]���uC#���3�`���U����j;&�Pf`�g�W���?�y)��9��8��l�4��H��D-H�'\��qK�o&�*��h`�l�4��H��D-H�'\��������?v"n<�#Ƥ���y�I���F��*OʧI�8��_/N�c�{�ty���
�<��^�:�)_\���L>�~��:c�gM�,`���<Wԭ	ƽ��~wD[����B<:����t���
5���4�~wD[����B<:��O������p.�����4���Z�u%��;��x��<�����`B�)續\������kD24�ͻs�	Õ�)X�JK�IE��́	P6���4�ͻs�	Õ�)X�J�&kx�|���W`���?�fpx��Pp�}��
KgqZ� ��ڧZ��7 bt$}΃�?�o>��!`�u�!j́	P6����|��{�r�\	��rR�{_�3'�X�)��}�OVB>l�2������[u@�59���_��ƊH~��j.o�c�\.U1+]���]`�Ү���3t4l9�F��g,�5�TzS�@/{�&�_��ƊH~��j.o��)����n��3;�í��>x��F�\��Ɲ&��&0��n�~��j.o�c�\.U1+]�Ȯ��ߊ�X�� ������Rm�Ƈ��ݱk4# �
)����:�u�J�/kz7�Y$��S�*���X:�*��ܟ���"�hUioέ���K�IE��\���L>��|�%����0�3p,��ǈ8V\*�����7!h���X ��L�m�M������k���t^ꦤ0�7��65�Su����P������!`�"�X����GG�8��F��@���j`�;�_�2��B�>K��t��<�k{����Sc��6���y�=k^ŧMF��@������׋4>&:��Op��)ɲߵP�L�m�M����׋4>&:��Op�!�6l�v2�E� o��*�2>�1$��_w���<�Ú	P6����G�W�̩c��@�)���8�Z��|�����r���aM"���﹈�iklm�"&������r���aM"����y�j\��3"��0�;e5V�]C��%��Ob\���L>�B%���O-�#���[�?�c�	@x���1�|�c��1��;b��1�)S��#)J���l���\�M�u#RRklm�"&������r���aM"��^��J�Y�y��{W(3���P�^���������r���aM"��L�U���;��n�^-.�T��s~�U j=�	"����;e5V�]C��ؽMBW°��P'Q^|v���Q�cel��oW���3"��0�;e5V�]C���[���?S�*���X:�*��ܟ�tN$W�ٯ~�PJ):B%���O-�#���[�"yd��N�}�g,�5�TzS�@/{�&k���<9*�U�C��z��-p�Jj}Ѯ�/ښ[Tklm�"&������r���aM"�������4�D�Gۥ������F���9�@Zd��`�H�s�# ;���!��ZB��,�Ӏ(�ٜ�U�n~qbS�xǠ�j�|�K�U�z��e�K��2��9�냂s��Ę�}��U���)���w^J�b�=�P��/�f������o�rA��$#J7l�"b��"Z���RT���ڋ8M�.�<���Xz���0 ����o��:<�w�xF�!���Fi����oz�g��� L���dL7A�k�6�Ѐ���l+sj�yIZ8M�.�<���y3�/q��5P^�\8	ĕܵq}f=s@�&eVC�8M�.�<��Hސ��e;7A�k�6���BL��=!�bZ��b�Be��ڡ7oA!�䀯�5M�G"�ˏ8[$0���&�nP{5��_ۑ;���A�Cm��b'&�3hǴ�� #��L��_�wb�md����*��Z����˴J��sr�l�q_����j��?��9)����`\F#[X����[�B �n�6ӌ�IۏF��Aɛ�(�P���9T���l��j���^�B �n�6ӌ�Iۏ�+��G��L�K�=\rۤG�#r�\���(.�"�_�Ƴd�����ca�\ź�G�;e�|����p^���N�����.�WDv�b��h�Ӆ��x�����
�?<J�!�Ӑ����mi�b�md��/����h#Ȑ��t���13�3����*��B��������:���N3!�o�{�[�$<��D�V��\�W�EC�mg	}��h�6Q�7�y["�W�����Q�S^��c-(���mg	}�	W��^$k��]I�9�\U2�~xao!f�	�Ĳb�M� �{n�UYڕfC�(��EZ 4b�zvѓ�w7y�j>��l?
�A��t��#2��S���^RSŞ�Ӣ����NǄ��^�h5����N�U�/r�B�,{�d�����ca�5�B�V�)s[�3��kd��p'k��o��`��[A+��F�ڪ���B�4����0��GZ��-&��ح(��? "a��.,��G���B �n�6ӌ�Iۏ'�TI�A��8���9�GKP�2�����Vc2�����Vcl��w&� ��O�A.��T���p��h�ocF���(ZH4~��2�����Vc2�����Vcv�iL�DLV�4�ұ��ݣW�]1?�g��V�$�r����[�$��������>���3 ��������n�Z��b,ܾ$�m�s�>CCMyo=eK��G���^�o�A��P~��_k:y8Cg�'�Z��b,,r�%*Z������G��C�0P�@��*�|lC�r������_��}����4�]��Z��͟��`Q�u��E�M*G$�ץW��xl��2g���z`Ε�ھ�i�䰥�R<\љ���0e�P������&T�ͪ͌nU�B%7��U�ʳ�$D����s;�z��E�@ ���:��`���g<�:t3d=�C(���Ty}�"����q������_���V'�g�P��t��N���*UV��o��|1��.ٴS��@K7Td� �*ZJ
(�� 6U��o��f��[���m���ccΝ���0f�M����-�f���meD�@����-f#8�=��=�I��0f�M����]v���ۙ���-!��0�,W�T�!��c��>,���*J��L�]�|/g�����;��qV�F���AU Y/��'�Sl�{x�m	����ԑ�M�
q���nDJ�t���7�ۀ���3M��B2�k��u��t�y'��BS�5S�7��M���5^s�a�O��[G����Q�?ë<%��KM�!5P8H��E�7/ �˅��B�,�%�	w���.W�~�����Q������9��̵���cJ�ҽ�V�hV4��W˝�ѷ�[�t�V�M���5^s\��M���	�k�gQuON,./�����o�����5S�7�X:[܀O1�ԠֱTU�49�5�{��8Y��潇\�k2A	�\�t���a�A�Wӫ<��\x����i1��s�$����ns)��E�$*:e1�[�"zz��T�4}ݫ��%7���� ��#��� �X֐�K�ҡ�v����o�����s\�)"ߌ���F���֦V][�����yoZ�P/=L�X�s�� ����7�ȕ[��f�o~����RLT��=��R���3b�����d(P��<��lDsN����p\ט~��Vz��lMV��*��o30�@C��ǲ��7�{�F�T�xx���|��*!��	�6�V�Q��4�d��Au�{�|5"E&��� ��l$����
Ő�G:!V��,�O�!\�"�X[{�2�L���h��N�U��W�*<λ���2%0���#�͍�rko�D��=�C%��
|�5
\-��Y;��i]>F�����Z��+�d}ꑱؤ}�Cğ3;5��}�?�"3�3��gL�G}%KkkP�ǴB6²7>��υ2�2JTC�X �� WR	���Kէ�[�Ǐ�9���)
��"E&��� ��F���֦V�!n����sۅ�LT�(n�l����8�^.�ܾ����Ҧ��D��ܒ_&^�� �$�^&���.����V�� ������h{�Ӫꬕ���ľ�OX��ʹ���r�vK;�Af]^�����/�@�h�v�9:�8��yg�%��=rFq]��V7v�鍾.�{C@o��@�rbt�k	����-L7��uC6��� 4�����0e��H�\��C��E�3�S�ϒ�eƀ�F�m��pRO:�'Mcö]-�{�����k۽!M��2�=�-�f���m��bK ��&Y��V�Ձ,���K�C"׶�Z�+՘#ZZ�sȸ�"rR��L�䎼�����
�?<���ilg��-8c�i�� ���>w�V�RDFR7�U5�p�+,��C1���(�ѕ��J��<�..�4��˺�ʘ�p���ʘ��=���"���]�U��5s���Z��	��h �7w��WN�d7%�B�&��Ź|�Ǫ�"9EDK4��m0�� �d�Hc���[=d<�V�QK�}�ݓ���;5��i��_.j��ۖ���3Y����� �k[�d�bș;��<�V�QK�}I�I�� n�6~ [�W�A�ޞ�ݮ3��������Uc��@q�;��g�dr�jf'E��"�4�x����-���[(P�S[W���w���9�m��
�j<�p{��{�-�RؼӤx�a^?������K�XQ��3����]���u��A����l����4�n���xǊ���,��i G��ΜޅKf��"����H%����e�r^�G��-^/��iIK��ަ1����rap,��~^�c�.[K��m�� C��+(���ʦ�G��m'K6�o8:4�p8,3s"=k�Rm���0��� F*,ƌN�jK�I�q����U�a�<��g�d��Z5W�
�5�w��L9��|,��[��D��ܳ�J�ʵC<�#�����o�K���d7Ud���Pn<���#�K4��[Q���d7Ud�S�CП�u�>����9�U2�J�D��������d��K���<�O�f
��y�J�#z�P�!�c�!�}�"AmZJM���`�D3��~��6��۟<y�׀%\N��qs�������I���5G%{�e����8C�8�����h=G%{�e�WOF;�Z�AJ��w���*���d��4D���tY=[�����ح(����C1zh=s�(:G��AJ��w���*���d����C1zh�Y�#�{U�x(�i��/R�������	սL��$Ó�[���2�����Vc2�����Vc2�����Vc�cRq>hb%�k]�s��w����KF�s�d��>�<^&!!HY��f��I�2�����Vc2�����Vc2�����Vc2�����Vc_ސ����q���:�!���p^���7�Y�Z����Օ�l$P�ĝ�ꏛ{{'oL�F�!���Fi����o�ޓ��-�!��Tӧ~�Q6vmI/5(Q�g�+%f���at�)��d��X��WG ���25t����M@3%��H��	W�UT̈́<@��L���dL7A�k�6��I�ߋ�-M�O��~��N}�}�����ߺ2����E����e��Q`���I\CZ]������E��׏�����Mx(�i��/R�������	սL��$P�V{�]И���
�d�����ca�؞�����L�m�M����׋4>&:��Op�������� _��s�֙f����h�Ӭ��SG�d�����ca�3*>ۻv�!wye|� f�Lu�m.w[vB�0�&O�;u��M��7{��(:/�b�&�q��ax��Y�L��x:A4bI�s�U�q �~k�%��x{^4��*m�D�$0��X$�����gtv(�Va�ir	W��^$k���P���g�d�*s���j��։�s/�V�kam��V�RDFR7�`h2#25g�[䅚˞��\�G������A��׋)тΪ*�V�Q���a-6�Da����
�?<v�U����CB3���K�d�����ca�3*>ۻv�4�ڈt׏�����MJ�1���۪	�}a4�������3'�L�N��V_�1�gd*�eƀ�F�iF��&��	W��^$k��������Zw�ʘ�� �hQ4�0x_�EF��sd�����ca�3*>ۻv�^@��=�6j�"HsA:D�D�6I\�zl��։�s/�M����� &'�����7y��c-(��l���@��8�z�-���4&ݞ9��h�xm��.�3���l���0�0�h��#g�k��g?	��o/���6��I\CZ]���UMc)Z�'�E�Jg�%o�w�X$���[�����NH�Ui"��B� ��~���4M̍����Q6vmI/5(Q�g�+%f���at�)��d��X��WG �����U��eƀ�F��*CB��k9Ӣ�p�)��b܉�����P���g�d�*s���j��։�s/�V�kam��V�RDFR7�`h2#25g�[䅚˞��\�G������A��׋)тΪ*�V�Q���a-6�Da����
�?<v�U����CB3���K�d�����ca�3*>ۻv�4�ڈt׏�����MJ�1���۪	�}a4�������3'�L�N��V_�1�gd*�eƀ�F�iF��&���h�6Q�7���yoZ�P/���ؑ3��^�h5��0����_I�����
�?<l
b���1*�R3�N����,�ǰR{~g�O"Z�#��������
�?<`��Đ1d��։�s/�e�*[�9��d�����ca�C�U2�����Vc2�����Vc2�����Vc��;����KW�*�	S,�d;vt����g: k��2�����Vc2�����Vc͞����C��m֐������e�  �.4^�&��t&��j�қjI�"��)�l�+4�]ed��{�b�IȀp/x��,Q��	}QorǟD�ui9�f?Y�OV�W|�B�I:׷�F׫�J��l� �[��׍��������֡�\�<7�X�e����]��m�n������"���P�`m��';��?2^�9<o�nïi��n�5�F�^hq��:�����Lh�7�Qa�_�G��Ǵ	P6����|��{�r�\	��rR���k�V�\���e�Q8-�^\́	P6���o�${U��w�X�|0��ѓ�s���O��['���x��U8��\���L>����e�� ������#��r������r���aM"����E֤�*�5�ٻ1�RR�,�*Ǚ62�3�����g�m>�`^����S,د�p�L������� ���8�%e��ڡ7oA!�䀯�8{+��
uj�����O�D}�����ņ�a�t��A0n���J��x��uqq9/�)�ԙ�.������Xuε�!>��/�����j"^�����ϖ [@wP=�	�:˳0ʓY+���_D�Q�C���� �
±2��h�6Q�7�0ʓY+��g�$��b܉����]I�9�\5">�E �9���=���˵k�^�pfn�R�k�ew���m�Z��-&�-�5�H�^�i�ӎL*$c�\�^>ZObW�!�
����
kX��!��ೣd5�͐��%�v�x�zIb�E�0W�l�l���XU(�a�+93��CxO�`
�-��d5�͐�-��;���:�n:G�j�jz+ ^,e(}�S�����4�֧��L_Q�����f;��V��m�;Ź��'�?�j}�˵k�^�p����X� �Sy�A-,�:���N3!�J5^�ұ�|��d��w��L9�ۘ��ҧ�?�\���3cx���K*Fg��,��˛AHCO�i�?��kR�KB��}�)�<��D�V�}Q4XʰS'F��-�x�h�6Q�7��m0n��,�0�wg%c�ִ��#"�w�Xb<���h�6Q�7�2�����0/zﴚ�:�L��?�<O���e�|���Dsw��J�����:��!$��;�s�*�:�L��?�<O�����+�	����X��֑xGVָ]���=A�%&^�nƒg�|R��qMw�}g��ti4c�St��'�r��'q#�� �[N0N�b� 0e[O��ɔ�<5���3g6�9
��G���1j|g[Ҡ(Y�u�/r��#�<���=��s��Q>�^2�����Vc2�����Vc�Z3߯���oL��ɭ�����Ni���2�2�����Vc2�����Vc�cRq>h�a�{K���6B\n���Ϩ���]k�kIY��oBd?\$��M��ݺ|��W�����ώM:��2�n�ڤ���[U�&�nЮ��\�]\���e�Q�����k�/U���!-�iP��G��\OL^��>%�Нo@���;1?�[F�9��G:([9��qUB������Wi�g���h���R���ɢ���ڠ�Q;�m��j"^�����ϖ [@wPcIn-Hzn�!��ZBV�RDFR7��D�
p���kg>�[OF�ѿa@��h���R�޶(xʶ���H3=-��7��k�VX��he�	q�X�Z-�_���mA�N�\:����v·��E;�ٺ6�w�н'�o�t��;��"h#�)��*N/�p��>E��ѸZ�����=[����ѵ�������?��ًGx�6��*B4��c	�yE�,�I��ގ	�� �\|��Ea+a�G3�u]˴�����x_��s�֙Q;��؆JWJ��w BM��ɋ���C������]��<a�9g�M�G�nE�̜��W����u�u�d!j�e{�~��j.o�ѱ}����S�U<f9^6To�${U��w�X�|0���ߪ��w�����蜗��,�ǰƺ��kÄH_��#��aѤ}[WckL(�Y��1v2��W
_F@SЙ� "̧�Y��\|��Ea+a�G3�u]+�u�G�k_��s�֙Q;��؆JWJ��w BM��ɋ���C������]��<a�9g�M�G�nE�̜��W����u�uPs_*�GqW�w��fD/����p���_V�r��%��;�tI�g?	��o���Y�]~p <�r�\���U(E�pOd<N�!�Q�f�:3b��J�Ve
�AOWm;���:Y3Iz�SŞ�Ӣ�F��������Srٌ�y��Kᷪl?
�A�� L#_/�e-M�O��~�y�J�#z�3W�ǡ¶֢��s�Kȏ���*�o!f�	�Ĳ� {�'#��T۳�͕��AKd��y c�gtb4�^���F�f�J�Z�G�O�(J��w BM��ɋ���C�����Ӌ�T"��D�x(�i��/R�������	սL��$���7'���I`����%�XDH�tt��ig}@��Q��)I��B��7c�p�V �!8�8C��z�:Y�����gڟ4���I`��y�<zQ���n��뾦��c�������C��#��>��:�@U�g�q��}.�WyT �$:�#��>��:�@U�g�B QU�Ka@��Q��)I��B��7c�p�V �pf�� i/�={"��sZ���Y�!�#��>�a$�i����c�Z�~����,�ǰ&k������ǆ8�ҁ��Tŵ�$R�i�Yl-)@xz�:e����
�?<.���6 �pN��r��<Н=.��E�E��Z�2�����Vc2�����Vc2�����Vc��Y7╙f��/(ޮT2V����uV(1тQ���3�u�l2�����Vc2�����Vc2�����Vc��`���4"�A^�F��gVE��Qx�B��������e���F�Z1��}ٲlY�T5�����=tQM�_����6��LM�<�>u��N�x��e��k�7ܬX�"�Hb^�G�𿫺}Z35�V_��s�֙C�T&L�P e�mC`���j��k{���e�V�{��$���G�"�M��.!y�O�|�5�<�..�4��\tb�Q��b�:�	$?�����e�>64[`�)6��9��xx�rDc��/�;���)�v������t^���\�}]C^�5Q��R���|�ޣ�W�]eeݐ���м{�%GuN����A@�e���?ͧ,�EXt�|p.�����4���ZU.⭾)6��9�ߺ����T�2V�q�Y�;�
��+�d��[{���_,�c$�N�1E��Zi�DЫ�5�|���XԦ,\ަ�It}�0�.�,��.0b��V�����c�,�%Dv�y �谝��X�e��}�g�{wln������Y�
� T[��m��U}�	�(��Q|3�r�^K������О.�!H6F�� .�/'�b���' /��~�;����ɝ\�!2A����ed���M��7�vsi����WG��6`Bmy;;���0��0��}���'/e����'3Ȉ�7�u��\<g�
7�����D�nR�����,�ǰN����;��Y߸I~H�1u$���B�����(�m��w��l�U�C��z��
������y��ٓA��E��锏��Z��E�ㄪ���wM-X����痴�y��������z�	q�JaQ�Hu����i&�L4⭦�����.ƶ�~b�!j�m�.��H�$��=��$�R�nl�;�w���vKz��+�c�����|�\;͖�kYIį�a�y{�הr�R_ǌ��g�0�u\=�~ o8�1�R�*���M�,������3~I/��\]��j�/A=�� ��u��ۥ<ab�۹��{q�J��pc,<�,��
��]�/HT�Y�[V��M*�x��<�����`B�)續\����'ò�������?��Q�&{��8�a�;"��PÛ˻Q�0+�kΐֈ&������A@�e���?ͧT��w�/�Zj����£�&|d������/��p�!���Ct�w#��@Ż�&ǥ��a���F߸��S�Ȍ��	k���կP�*l #^��|�37�˱�5^7]fn�cՉ�����ɝ\�!2Aպ@n���4
�|��D:����[���F1x��7cd1�RR�,�*Ǚ62�e�zj'qmf.��X���/�nxL�J����/D�;���O�a\Y�����y�j\�U��\�7��h�ř��ޔ�o���y���@	Q%����������r���aM"��r�F�*�_�JH�q���P�ꡘYᔿT�3���oDU �?�o>��:C�?p{^�S�$�0��&&ĕ^$&�3;:�]��r���Q�q>x�N�$�=��e��$��C/��~4�K���a��mY��AKE�2�n����=�~gJ^&�]�;~�/&$��8_9`f����K �_"p���4~1��0�RQ�� og�6�G�8�?�Y0�
��G~�T8=̓x�R8D�}���5ܺ��K��ѻ�G~�T8=̓x�R8D�}���5ArɃ�_K�ņ�}h$���n�۪eﳉ̷J)6Fx@�]�����͑����5�8Cl8R�j\�/��ɘ �V�	��`��e�>��y^Ii��Ns��*��]���\OL^��>%��;�줦i�FkmG'w����������\_ks	�d	c�b�xe�s8A�iT�v��K���qE���$y̮��@e�2�$ߣ�g��~�4�"4D�/�k�_�|��M��VwF?�d�)6Fx@�]�r�I���\OL^��>%��;�줦WѶ
�3��@hG����\_ks	�{��$&XT������WѶ
�3��-�L��t�V���4�i��F�e�ق"Ҡ���>�SS�]�)����;\0�RQ�� og�6�G�8a�+�wViC�mr�,'�0�RQ�� og�6�G�8��g��~�	�7���&��d��:n���+������gyE�O��nie\OL^��>%�eﳉ̷J)6Fx@�]���������;�5�8Cl8R�j\�/��ɘ �V�	�-�B�Q0��y^Ii�E�A�#���ܰ4$b�q���`��%��*��b�&z|X�L-�.n*R,u@G��5�1;Szߧ�U4���&l@���f�sR5�Aw65�+V��@��s�1]}��Ԡ��T=�h5S��k[�=Uì�J勓�]�Y)����%���I����d=}b�T�x���hAE3�%�\Y�
Q`?�+G�	x��?,~|s���q�˼?"cQ�GݔO#�Z/��v
���쨳\�J�n厩�q�*�[#�P���1�gv��X���Ȟ��_�7��q��*���İ�Ewk}i��Y��Q��g��!��ZB]C^�5Q��R���|���@n�+�xG�3��	R'�6M��Hz.C���~����Z۳
0.��5�ź^����f�Z�
��>iXqP.W�my�'�r��'qm�±��m|7�7y�]��v�-c;��5����L���׼��8�4��Q>�x)��k\�7Do$�YY�6M��Hz#mԃw��#�r��8� �������iA'R�	���׼���Y�����Y'b�'=�(q��S%�d��3��4�Ef�`=�ح(��� ����hA���B.K�o�Od�"F���׼��]|��ť��z%�ژ�(L5ӥ���v��/���@�Wu�t��o�F�\���e�Q��	�2�R���Z��1S����k����O�}ZS\�n�ï��)Fa��V�x�l��1/Ax��}*���AUi@=���b���3~3�p#H*W��u�a�$Zچ��<b�Xϋ?@h���X �(��%�*ҕ/s7gX?�ᒹ�G�h���X ��Dxj��U�m��KBʞ�j�� "�?�:4L� S��/s7gX�.��Ԕ��a�-AK��«��N�%U�S�t�Z�#�j��1Lv�3`��w�E�V{��M{�l�v�A?Љ'�-0óWy������U�I�����hy�(2�q�ۢ�\OL^��>%��<�q�Y����Z�Z�\�I�\�\OL^��>%�P�^/�h�SL@�>#}�[������V��e�LtW��e���d�tAAI�O����09�	$}t�c{DJX</��G����>�]��*�?��CG�B a�޶�oo=S�
J1!��]c�ꃤ)7��lI�q{��*�5�ٻ�ڧZ��7H���hVJ������b	h���X �LOi�xg�|��Q;��I��y�j\˪�,Z<9V����ft�Ag
���y^Ii�qpըt����X����\OL^��>%��<�q�Y�.���x�D ML:�\OL^��>%2�C
d���Xm�NR��J^L���� "�?�:4L� S��/s7gX��R��G7�Ԧéc�Q�ټ:��N�%U�m{ xW�Ĥ�Y7�Z�����T��q���j���v���N ��Ʒ�$��+�7�ͭ�s������Y=��~<6���m1��%5K������L��S-��S��HY�V��"�Q(���v·���Vem.��R.p���Ԩ�*������:�ؐE@>���J)i�r�X����9J*]#IH3���ME�o;�琾BT��K�}i�e]y]�g��xI]�-����q{�X5KY%��ִ��#"����]���&�n�Bk��迿��!Sq�#�-��>�C�~�)`� ��q��._(��n�Y?v�<Sq�#�-�����ؾlSw��,;7�?�<O��� ��Z�!3��\(FK��WdM4@ȳ$hI�+yX>�S�L��ƴq�������L�Y&U%����f���5�ź���ɝՄ`��G�Ȧj��`�e�%R�t%>^����_��Ǹuz�4�+��t,u:�@�Wu�t��o�F�\���e�Q�������r���Z��W��Ws��>�C�~�'Vp��U��H�Nb�*Z鎬�������(����ﵠX���G�Ȧj�B�ek�5Wt,u:�6?*e��;O�Ҡ�"�tѭ��xق�������(F���14��������b�-W��4 s�#����"���f��E���#mԃw����YNg��?v���cc�u��m,3�y9v7������Vem.��R.p�ǩ��0{5�ck�Bɉ���o
�a�JU%����f���'|F9g�M�G�nY�cR~�/��S�aE�@�N�	y���m鵗p���x��Q>�^2�����Vc2�����Vc2�����Vc�Z�D�U�3�P;9�H�.	O�F��1�9�GKP�2�����Vc2�����Vc.�
͹U��@A�"Lx����(�"�4����i,ih���64R�����ޙ��] ,?IY%�!�#g�k����V9�C^=.,����k��˔�#M6s���f��5�P3 C�0Q���g���6�����x�l��1i�t�Uq�_���13�׍����V��ÑR HjlU5oܛ�	���G�˹Ď��'�3�$ �#^�Vn�����'MRmHX���y�XZ@po\sQQF�;�?2^�9<o�nïi��n�5�F�^hq��:�����/�OP�I^���V� D\���L>����������f5�%{��t^ꦤn�da*;�?��CG2��6_�-N6��`���ם�F�e�n�a\Y����_�G��Gӌ���dֆ[�$��X�aM0��x9@l���v�&E��t�)�8	�p���3Ns:r�vbH?ߐN���k�N�� �\	��rR���f��2Rߤ��:��*�I����(����Iۣ<�;��O��8��͘�����9���F1x��7cd1�RR�,�*Ǚ62�e�zj'qmf.��X���/�fpx��`V-u9�`�klm�"&�&3�-��_ih�7���ӳ�Y�
����.C���SS����� �GQ��i=���[����)�y����|�u�{�غŋ��6?L��\���L>����EW����:�?��y�j\�ʷ��&3�-��_�,�]��Κ�3�ol�+�\�p!|T����l��;�4~���;A����z��ߩJ�9�h���X �Z�^6���t�Wq��iQ<]�I�ڼ<J-Y���".7�4F��(��z�+��p�,�#�w{:IxoҢbu�ߞ�(ɡ��'ƌF��\�)�`"8M�.�<��7 9>�B�u��m,3ĕܵq}f=M�C:4�ָ����Ɇa����:�;��NXv�BX�C����Q�_�N�g���"<���s��]b�$�Qen��M@3%������#�Lq���Bl$P�ĝ��D����z/5�L?��Vf����aUZ���RT�����h=�R��a:߻�%�q�i��¹ ^��y}$�)`� ��q���iZtO��F'ot#�r��8�M(]�-	��\(FK����HEc*3���}���Y�����Y'b�'=�(�#xJzc��*���d������O�]���=A�w�����a����gW��_K��Sq�#�-��� œ�Ę�:�n:G���f�2���7�9���������D�iF]��v|�ˑ����p|3��'�)n�J��N}�}����1�G�Qc�k]m���~�ch�Gé�ĻP�q����W�7J�Ka!s"֛
.C���~���J������H&X�J���o3c�-��;���:�n:G�d�4�t��Է'�r��'q#�� �[N0L*$n�
S�}r�HDʞ�sB�_қ^㒤�"_��Q�$G?����,�ǰH7"LTft��c�}�!����ޗ`��K	���o�e/b c������*������9?�d���&�M\R�'��5D��0h\Ef�>�"ª���Ps_*�Gq�p���x��Q>�^2�����Vc2�����Vc2�����VcEb뾯�J�UF����0�e��#�[����9�GKP�2�����Vc2�����Vcv�iL�D*M
�Y�cY��K�^ �)G�J�cbp��'@
9��y��%��3��׍K��ֻU:�BIWu��T!���I�Y��Q�9؜�%�FM�'7sNH�i2Kq��ٗ9؜�%�FM�'7sNH	@p-��Q�]��TM���K�+EC�A�w�(�XVb�w0[�؋��ګۗ9؜�%�%=⬚��dhil�C�����/*8��������hil�C�����/*8��״�њ���zͳJ���%:�q�������
�):
TTTW�Q;�im���M:��2�@���U@���:��F���Ed8���d&(C�#�7#^�Vng�m>�`^����S,�X�*�7>����p�*_�j���V�2��Χ�0_2b�� �.f�8>fd��#��rݮ�d�3a��Qj�[_�}��GN�`��B�0w��zw�r�Y��nf|FN�7�gI����I�}jA@}(���V�6c	�	r�������կ�>	F^����h4c뵆qR�R��Q���J���3c�o�����h4c�Ү@;���!��R"@�j���V�2sQ頭q�a�t��0���v`�2�����Vc2�����Vc2�����Vc��Y7�8���O�T�J�UF���0�C��Z*i2�����VcN�1�� ��2�����Vc2�����Vc2�����Vc�ׇ�xX���Vem.���9!h�V^�"
�	��dvl��?���x�l��1y���ri��nU��X|Qeu��<�́	P6����G�W�̩c��@��O���l`V)�l֐�N�T!ߤ��:��*�I�ͱ�U�Lĕp�fpx����(���M��oP�8��e�*���|��t��\nq��4�ca�(f����j�ơ9��&@�E�Ws�!R��p߷Td��#��>�(}%@��7�����Sq�#�-������&�eq��˪��c}��-h���X ��Bw`7����w�Q���Jg�C>�h���X �i�S�E͂��Dc�!vj��dǑ؆�!��ZB4���j��e�	q�X�Z-�_���mAR6�.�iGJ������y3�/q��f��n���t����K����r�5+1���K���<�܏�1�\�s[O��ɔ�<5���3���;�W��녕@�E�(�����6N�T�f�'�r��'q2I����J���T�D��1�G�Qc�I����4��l���8۴�k�8v����]��s��/� N��r*`�̮0w_F��e�������ӡ�6F�!���Fi����o˰]I��x��n�bdk����bup���V�[3�.C���~����Z۳
0.x'�M�h$��1�G�Qc�I����$-v�Ҧ�B��u�u�u[�z���IX4���1j|g[Ҡ(Y�u���LI�֗M��EכPT922m�F�	�a2(�!�f�hG y�7�[�`kr��&R;V�
�#:�L����R�����gVE��G%{�e�WOF;�Z��I 0�V���bU__����;�N:?y�gc̖�)�p��6����Y�-�_{sx�L�}B>�u:Q��v4����e����)xZ
��+�8������^{����zc�K��>R��o,���c�K��>R�q�Vٓ��(�����ꛓ�]ɞ(:�����Og?6����V����J�����Bw`7��#{63�~}N�cPb�D�5P^�\8	��c��
�l$P�ĝ�� �����%����*�E��M@3%���n� �Q� �:W��Z��Og?6��J�
�Mɷ:���N3!	 �����b��8˛AHCO�i�?��kR�K=s�(:G��o��"���h�6Q�7�
3K������&��S�)��X^�uw�c��l�,j�D�?_�3˭���߈�vJVt�l�褻�sv�Ο��sP�;��|Bo'�]��ɹG���Ĩ�_�#��� h�",oMG~�4���Z����Cf<s0+�pΡf9��`�D3���Z�/�0��)�P؎ߤ���&�E��"+VqS?�d���&�~S���v���G�����l÷{H�D�U\���<��ɄQ_���'�8S�E��NJ/��!�#��W+Δ}M��R����0�0�h��#g�k���u5�E���9I7�=?���L�Y&�!��;�����L�Y&U%����f���5�ź�IM�P�Eݽ�"�{��,�ǰTm�v��G�U\���<����${���#'26�-M��{w[�2�����Vc2�����Vc2�����Vc2�����Vc�i��������J��yԴpZJ\G!@)c���Fu)n2�����Vc2�����Vc2�����Vc.�
͹U�pϣ�و�y�ݱ<s�n���s�w �9�"�GC�N~,
e�<�V�QK�}�j:���`+��~'2?�EQL�������D��ܒ:�5t�W��{%hPb�|�������QB�'�KW@�=�:����5���֡�&Y��V���O���:��o����3�MD�ew�P��Xu(�=]ݮV̆s-Z����Ѯ��l���sGJL
������xKI�� �LfE��!�&�k:����R".�����''µ,J�l�/�'����&�"�o��o���Y�T���6��3m�G\(~%���=���[�ك��N̹�Y�PG�(�Fn{��J��[�n��g��\Y�7�
Ύ����'��%�v��6
RS�8���$8�%���./4q��M�$)'��:�Jl]N
��FmE�S�h�� �Ѡ�˰�O���:FY�_����c9S��D�j���r���I;�śE30�A�zc��i����T<��y��3�-N]�����$h��܍ˢOh3bU��*����b�[�Ҳ۩u_�d����*#�IQ܋�w�
�`BB$�W%�@���&�6L�'�1DcЌ*�@�c�.[K��m)�Ty�cR?�����_�zw��Mٌ�ؔL�F�W��	]�	���D��ܒ�0�Ex��_�j�H�#�Q2`��q4E%p*�7�)=�zxh�	�bC�/pfNw�&�Θ�xw�<2%��O�@י�m4�1�]��e���im���2?��.?��	�Ï�=7�}|��	D��X�*��_?�v��9�2�L%J�bb��|;�����8������t���MIV��8Y��I/��\]�3�� �frw�ܲ��}([��}qn
V~$���ȏ��F�[�c�Ĭ	�g����#k�˟ܒ�o|k�Lb�5ߧE4��J�1���k_���b_!2�͞nOYԐ���8�H�?�#�=7l�"b��"�c�<��uS�4q�
��?t�+)�t���(�x�@�
�����jR&l���7A�k�6���gݸ�$i�����&�½0�M��h�6Q�7��^Dv�H3=-��7�,
��0B����/^�À<MN2��΢NE���������=�T��"�&�kc�
^	8�Y�&�jW� �瑴�rY�g�0�uk¨�Γ�7A�k�6��I�ߋ�X��WG ���zt��[�h�6Q�7��^Dv�H3=-��7��[��9�΍�$pt���t���(�x����o<���H��m�Ƞf�����I A6˃rG��n|,�Rn
V~$0�%t$jp��v|�ˑ����p|3�o}����ĳ�e��@N���Р6�#�fp�J�ð��T��~JFNǭ	.3y_�r����0�E>��\9�oA$'�J��>�����&o�γ�hI/��\]��rX�;2����9aP�&�kc�o}����ĳT۳�͕���zt��[�A�qL2�cU�:��(�J�1���k_���b_!2�͞nOY��Q>�^2�����Vc2�����Vc2�����VcREBR�hHr�mi�=�ŧ�٘]E�)�(#�� !�hr���2�����Vc2�����Vc2�����Vc�cRq>hLV�4�ұ��but�;\�D�s�,��n�uȓ[������M�&ݫ��W6� ��\���<�(eGq�����r�����T'Vp��U� ���sX���4C"1v��'\�|^�^�h5�����H�.�����
�?<��Evt�I��b�F��x����X^� $)�lj�iE�EYZ/�VU�簦-�b�+�