��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�|�#A�)�(F�ow��M<r��`cbp��'����Q4�^v#ȐUD� �m�'�t�חEʭ�3�Jl\'q���v�/���m���B̑!<�!$�U6�b*��G�DRf_��]JO1?>����d�I�`e�D�ǖ]��!e����>�Av�^6�ˊ��Z�]Y��8z(���Fb����H��G4�"n��O�䓟�&ݏ��A�ꐖq"�\�4;�g@,+$\�M�h����*�J����{��� �l��^��Pʇ2��"Db�O��=i�Yr�a�n��W���b�����j��~����/^�wG$�Ѕ��M����W�8=�{j���g���o�e:�Y��J���F�H
���[F�!e����>j���g���/^r��`��w8=�S���s>.O�CSeu��<̎�ɤ��C#S+�nʥ1��9C�.�^<% ��^�e:��/j��Ψ��F�M��;˫5+J����T�)�[���<�L��͗���X�#zt�d�1�� 4>�[�y'�y�� �s��ɤ��C#�q�^���'��a�"��Q�u�U	S����o�|�K�W-��vu�TS�m���=,�4����Է}�š&�c��YGQe�.A�������ҧ`�2'2+q�z4�m״p^��gs�N���Z�0��m���Zz�20k?�i�cm0+�
�6�.�)����/	e%J�bb��||�G8?6��ת�/�)�I¿�l����4�����Mq��}/E�������ߎ�� �:���	�H���i��П�i�$��x��F�;�`W ic�ˉ-W��SL)��:|[%.�m�QA�Q* �#m�*b{��a��n�d*����l����4�e�kzP��cA*�["thv�x&(w{�3��0�أ�M:1�#���J��E�	��A;��T*Mv��%�����dN�<@Iv���a_|��������7o��v�3��OңJ�<��6�.�)����/	e��5�ͨd-f([��V�H��X��H���z{<���낌�c�Z�~���ŕث���j�)䔫�d*����l����42�W��x��xn��/������A�:y ��@�>=��}cbp��'��cA*���̟��cm0+�
��ߎ�� �:��ǝ�JJ ӏKg4	lr��e��9�j���B(QR���ScP"Nq컰5�&�z;cR� m�Nw^x�p�]`Cp�P���/R~dU&��(�VxM�T��}���.O��#)]��.�gP���n��8�U(���/�)�I¿�l����4�̎֍C���o� T���Ig`i��ߎ�� �:��r�Д� �}ɧt�A�{*�}���.O��#)]��.�gP�\'{�B�B�U(���/�)�I¿�l����4�n���xǊx2����0蹝�#%%��t&:���aKN�-cX��\'{�B�B{P�O�>dG��n;U���S���RU���Wi��L��#��|���kJ�@�>=��}cbp��'�+��^Vǽm^��`2dvϞx�p�]`Cp�P���/�%�i0�i!�[Oj8lr��e��9�j���B�<Vo�eon�_q*Z�Q�u�U	S����o���AC[_��{�mC�K��[MԲ����;/��Ҡ�@���p��v��Rb�ybq�I��(}�Y�T�x���ߎ�K�+EC�k�~Z�744��S���Q�����F��˷��7�C��zC@O6��r���k�'�<�p��Z۳
0.lr��e��9�j���B���M2�=쪆�h�L$b�M� �{�@�>=��}cbp��'Ӡ߳A��A��j �D*���H��gx޲{�ؽ^�>��6-k���P5���F|�MJH�K�{HLw�a���`�;�x�渽5�����z�����-�0ᯋ�q`�he����ӓ����J��@b$�(�1�M:��2�	����t�\�7P��T���˨�O��ܨ[�Ĩ��闇�:ۋM�7�	<f��&���x{�:AO����k�*ί��8Tˮ�o�9�����������ҿ:�c��k�?1�4��|9UN2F�찌�j���g��ǁ�*� ��1��_�y[�|�L�M����2�tj���g���o�e:�Y�NE���a�j��]X���{�ɱ<��5*f��.-�U�d�}6�=PH
���[F�!e����>j���g���/^r��`���HI�#�Yn�Bn�W���29a���Q�0��;�E�Ģp�ҫ��KALN����5�����uw ��iȎ�ɤ��C#�<��Ȃ�?BUY��E���q5�n�yG����y��Ψ��F�_N�瓗��ƾ�,oU�"�J���+�&�EX��K>�\�:��19TH��@!Z�p>L����B�﹈�iQ���n�O3���##��P��Q�K���F��ϓ�� MA�0�͗���X�#�Jo�ug�ZQ��#����TF2iг�Wv{{k]�B+���',fO�R���J1�/$���wW��SL)��:|[%.�m�QA�Q* �~�%yR͗I���Vܨ�C����摤ߎ�� �:���?�K8�1�~{pn˳Tlr��e��9�j���B�X7���w��3��u�!_
� �K\�����D�FUe��q�}O༠d*����l����4�e�kzP�
6�I��"(I6��f��Ig`i�6�.�)����/	e�Mv!���x��������=�\[LW��SL)�q�����f-��9�K�1�@hG����:F�X?��B����qe�@Rv���|z�ä�@�Z��&61������
_���֠d*����l����4�e�kzP�
6�I��"[A�,�OS?-#�� ��6�.�)����/	e�Mv!���x��n��8g^]c�؆�H��T�cbp��'�����U��G=X��������j�ӂsZe�/�)�I¿�l����4	Ve�Ew94�ċJ�obK�����W釵;/��Ҡ�@���p��D�FUe��q�cd4l���o��H"
��ߎ�� �:���#m�*b{w2���Ǿ�p�+�� ��	*vM�G9�j���B(���]*L��Id	�}�R��M�/�)�I¿�l����4	Ve�Ew94:��Ɗ�B<n�Y?v�<�;/��Ҡ�@���p��D�FUe��q�y~�oԎ}���.O��#)]��.�gP����M�2��R];t�n�?-#�� ȑ�ߎ�� �:���%�i0�i�l"����D��n;U���S���RU:1�#���J��E�	��A;��T*Mv��ޭ�;���Q�Y�F�
mG��ڋ^4"GKwHx�p�]`Cp�P���/Q�Y�F�
��6�ލ`��}���.O��#)]��.�gP�^��/c<�ja������n;U���S���RU��:?4sۼ�MT(_��w�g�P_���@�>=��}cbp��'Ӡ߳A��A����9��ڞ�7�2�"�&��3�(���e�&���6�$�5�ؼ��A�����x�p�]`Cp�P���/Q�Y�F�
q�I��(}�Y�T�x���ߎ�K�+EC�k�~Z�744��S���Q�����F��˷��7�C��zC@��)5!t�I~=s#�N��m���5�D�/�S���RU��:?4s�d�}�`���b�8*Dulr��e��9�j���B�<Vo�eo�T�c��TM��?\b����NfF;=|-�e�)��'���/(LI@Bc�~�1����g6:<��k��N�Lr���O]ݫ`����a0�m>�5tՓ���� }ikw�mc(N��5pd N^gp��s���+�� �#�pՍ7��q�?Q��c�z��	 ���O��S�7�_l�K��J����{��� �l��>w��;�W@k����cF��Cb�o5B�C�g�?��s��*o��^�w�r���	{�߳܎��Q)l��s���ߋW�(��?��CGj��]X��4��<L��H
���[F�!e����>fSeA��}�~x�K�0�F`)�\��@hG���﹈�i�~�Ԣ�s>.O�CS!U$Y��� ��dW^�:\��K"�NU��e>�5�����sGv�v�5+J����T�)�[��n�I�7.�rS�?h?���k@�����o��E1w�sO�?�DB�P�[1�c�
�0�e[�9�x��s�s!�N���:�|�z��J��
�@!Z�p>L����Bh�{V/5̏6���}Q�u�U	S����o�
�������S���Q�����F�π�-��pt`���(�ΜȠf'F�d������"�"7��v��� ���J�Ҝ1�}�R��M�)����`z�20k?�i`��e@�-�:�f�}���rfz��	;愵��Z͗I���V��T_c)$���}/Q��RU떐�ţ�CM�<L�Bza���	�H���i��П�i�F`����J�[��C�xMq)2�����H���)k<Q�Hǝ�J��|���kJ�����H�(I6��f�V��0q["thv�x&h���X �������S�a%�������
_������P��
��g%�l/�i�y��+����ŕث���a��n�����H�[A�,�OSsaN��@�8�6Dh��6ÈH^�\'+����ʄ�Č���J���!P�����A�:y ��8���R���6�ˋ�遙&�P5r7�^�~w���z\n9~��1}x|�±�3�����7oa,����gh���X ������'�c�������	��j��|{P�O�>dG�8��O�0j �L�?�A{�ا��݂t��] ?O��C�2�7��P��
��i�j9�򂃴��C,���n��8�U(�������H��nܶL���ŞU��.�]&��p�X�J�{��R?��6�������K���8Lg��1�R];t�n�/�@�g�Mc�>�W9���P"%��_��ɞ�-N��BD|�	�76�X:M2�T�I�]������C�yQ�p�E�U��
_���ֺ76�X:M2q]���K$�_���H�%�i0�i`eҝ2$�4�����L��#e]y]�gd�}�`�۫�j�)䔫�76�X:M2쪆�h�L$����)꼝MT(_��w�g�P_����aE�R=G��Aa���v��Rb�ybt��k�|�E�-�a����J�z�k��%�i0�i��DL:�KJ������d�}�`�۝$.Ë@�v��Rb�yb���<Q N��D4�ky���aE�R=Gm�E�)�J��!L#�]2v��Rb�yb��ۅ����t��#2�����:^2�	 Ⱃ�=d��F+r{�γ�5���$��PA!N�'�y�G