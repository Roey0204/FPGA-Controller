��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-?H)t� �hz2��ƿ� �lJE�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hp���Ť�Mn��X)r����#�L��P����⡇~g�C6҃�2Ee�Y�R2
�I.�%�$����o~C5R۱�JE�{�%�1�Y:&e���s�{_�1�1�NO�}w�3!�`�(i3�>=���#�Z=�į}�z��eU�4�h;��*�cT�� $"%�G�����C'�O�O�J�8�y�wⳘ=�C. ��f?��s^�xct��_Tҥ!�V��NR0�����O�,�WNT�N D|�5N��]V�'sH�{�����M�D���dle�oI�B<r��d���s�)��[�Pr� J&g~�������~�+��,/,N��$�H��t]�z�ؗ��6�����r�>>7�*�� �W9b�(^�#�s(Tl��d2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc&�ʖY��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc]�ԍ�[���S����Mg6�	�w��)�=���܏B��-b �|�ć�H� ����GO����H�x��3��O� ���&�*��*1�H�%����;H��F��1�+un���踩�#ä'AU�3t�R_�f֓�Ґ��1��Pld.]/t��L~�:��bۓ�Q$��J.�U���P��Y�����a������f�������n�A����&f������Ͽ/fE���ge�qZ��1����J���W��t�\/^�ɬc��WNF�o�F�w����?�<�V�QK�}�g�e1}� Ք=�� ƍ�ge�qZ\�h�8اN�<�>��L�0�(*�&!Yd�/�S&�z�E4O��nc���of��WA�?���m��G�$�+a1�Oj�ϡ����u��z� ��wg|!P���b6���Qy�V�SK���B�붋"�M~��a��J�'s��"|o	���=l"�,�>E��&�3�y�2��J�J�T�S1(_�'�&r�~,ptQ��k$Vʴ8�ta>!HԴ��ښ'��f���z��ÛK�lN��D��-SV1���A�G3�2��.A�_}��]���2z!5���sȸ�"rR!�`�(i3!�`�(i3UJD�P󹦜���R�8m�����-nԈ(��Y|	��7����e5�kFFu�ks�Fl�R�f�:��J�~�;�S��(�ze,e�-L��@X�h,#_S�3[�U{f�˰���&�3�nd(P��<����(\]�O!�`�(i3!�`�(i3!�`�(i3%��짐�Cq%��k�`�?��<��|"��[a&
�RY-�?�U<���!�`�(i3!�`�(i3!�`�(i3�o�,�,�Z�(��{���X�B�⸭�Y5p��`Z"�A끼�"�"�A%o{?��|T�#y6��
w� ���ѡE����mY�?�AO�]ׇӭ��!�`�(i3!�`�(i3fxkY�Eо��PW��\�����8�b��������!Q��X�e��*^ɍPbB0˩��K&3H2+l'�J���W&����ˋ7Ѵ� ��f.��3Y\c�@��#����U6P���GfX�>��JP,���[�c}�sXy�'�H�\����8N%�J�G��x�����)��ཡ��!�`�(i3!�`�(i3�ݓ�W���`��8Ykз��@��i`�T�Jp!!v*!����ܷ̔��aS�oAG���v�ͶN��B�c�|��0��aS�4��в}��aC�2V�V��"k@:GN��k�z���(8@ԅ�'���!�`�(i3!�`�(i3!�`�(i3��L��[Nh9�w��G!@)c�{�w�?�3K�<�Ņ�E�E��A�1pgx/Ҁ{�!�`�(i3�M�\�)Zw�C�'�"����e�cNơ�&Y��V��J8�����ۊ�d�Zn�T��@qsȸ�"rR!�`�(i3!�`�(i3�����hӠ����ه����ĜR37�@����v�c
�������Fnȟ�T��0IkT˱ �[r�vVˀ����)Y��ZU�	�!���w:��:B�9��aa�<^�>���o���o�^�d��d}BpI�ҽb��0�p�fb!��u�뫰v]uR�z��eU��*3M��t�[��(�2��o���o�"��8�O_BpI�ҽbi����ͺO҂�Z\iٽh�1{�/8'��taÓ�`�dz�'�u�Yb���$䀸~�W߁b!��u��\�W��mAUϕ���Ge*��]�[�����7��W`܈���hMo=�<*�֔��OW�6���o�� �C��I�"`
Iܩ{0)Vj�ꓑ2h�1�P}�jS]�רT5�'|w}�#��]�b��ގ�<>�T����o�� �C��I�"`
Iܩ{0)V���5�n�3����&�$`8�'�E��ZQ���޳{��K�O�n���(�S>���c��չ�=������)/(8�D2�j��rɏ��O���u�!��^JG�L�l����	\�R�&�-�"
길�����(�S0�4<+��80PS��J�aNSHk&��g�E�H7�81�Ÿr[�c}�sX�E-`b]�!�`�(i3!�`�(i3!�`�(i3���Jq��{��JVj%I��#fW�#7FEr�M���5^s�/�F�A@�����}���[N�)J��7)�c��@��5�L0gBnd?֙�꧀��*6��a��y�T��Z�Q����"�#&�1d��w��4܆XK�x��4����QXsw��؜�=��.A�_�N��2e��<�V�QK�}��{i�etK�y؄@�!�`�(i3!�`�(i3�4���i&�����^Z�Q����"�#�_.���w��4܆XK�x��4�oS++���x�{0��]�Ul���Βk�`�?��<ޖ�˞,c+�`��PZE�������!�`�(i3!�`�(i3�>=���#�/8'��vT����U�:�ƅf����V�p�_���ȃ~���'\/�(��\	wH��Y�� �k��^��Xz�	H4�����RN讍���V�m5�c@��I�����b2�{������7��U�:�ƅf����qC���6��������谶�� �"�R�-�c5f�/�F�A���_�Ұ�>��?2e��"�Na���VƳ��N|g�|��{�$�˽�Lk�`�?��<��t!I��w�d ��w��4܆��E�n�l�r�(e��b�αCg&=6�!s}6,�����{��6;%���;$��_���ȃ"4����uF�z�/��6�!s}6,�����{��6;t�|�AS��u��ߙ����Q��U����De�q/ه�����<�W.��[o�^��dH�M�$/�u��ߙ���¥+_�����|�Enz�<�]iO���<�W.�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����r���bW&g���&�V6\�> y2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)O��q$B����^Î�Vk��w/& �bRw�����IL�+�a�Wц�>��L��ʻR0�˧���.�E����F_���T�*'�uZ�ZQtg���&�V6\�> y2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯�^��N�&��?�2�1p���}������]�0�lK'���Xw��_
�u��>Oʉ�
Ү��p79�[vĄ4��5�������xv(�I��'�%9������kӱ�.��{�OF8�K�诧��FP��ߏt5<�
6�uE@��k����࠮R:;�L���9�D_�3���U_�+X���E9��*"v%)�(��(����������DGϴ�������開	����5J�^#9�<��\�v�w�?�b�>޼�\�v�GM
�-��y��5��f�,@Lo�l�8�fV��S���F�7Cg��-��1�C'��GW����1T�XS���`��Ƃ�$������cD ʯ6��9��ܰ�Hq�Ӯ>.��s��t]�%3������0|BH6A��fmO¶��r�``q��:{��� <&�M#�5y��;�;xI|$��YQ}P������	�̵<x
Ү��p7��@[��Y����J.h�+�*��C�����B��r���a���X� �r1� �V}$|~ïSup�xg쬉� }�����v鿪��U��ζ}̤��'n�^0o����y�] ��b�FP&
�c�,�%Ah�%4
>��XP���/e��I�]˅�UpQc\��f{u:~++��Z>H@��/l]�)D��*�V$ ��R8H�[��C��|�T/,wr�4�VĲ+%� ����������Ο2�K����3S4J�ϒ&�]�I�e��w��7;����#��3���Ct�w#��@N6�@P�q0M{����n
V~$L�
�k���۪	�}a��U�F]�pv�r���S}�>�~ez����開
���3q���"��yz,2�wÚU�	vn���D��/-�!ͪڕ6 �3RmRK��[��p^�g�O��̊�����a�"}�=Ll���՘W��.�r����m�q�pE�[xg}2A�/�����`z��V�g�0�uy
��Ϸ^�t(���k��?�C��k>?T�Nb_B� gF���D	��0�"�J�d��n�Vi��{C�{�2����-M�O��~��Z>H@�������1x(�i��/Rx��<������+�Ɵe���}�QU���B�ד*�h���&�E{������Hn[Y��S�n+��5�y��5��f�,@Lo�l�8�fV��S���F�7Cg��-��1�C'��GW����1T�XS���`��Ƃ�$����)Or�����5����`K��dx�b�W�6,;,塅߂�5-э����=���a֧z���>��RN#c�^iZi坝�=�G�XZ��QJG�?�y��h>7�*�,�t'����ş�z<Ҡ�"���p>7�*�֑^���s�Y���;�3"�Br�z�.�^s3���5��-��w��[�U� ���_Z�$=8�"��p�Ƕ�ڥF�NX��,�������|\%���=���a+��i�7k�+U�HJ�h�]�c���x�]�V��g� �x)f��p�b�z'hۉ)��Y�Z�#e���im�����<0�c��^�
E��4I-��>�!4P֡NPo��$V�a�G	)-M�O��~�+]�N/�|m���-FxV&,;�2{ �h�焩Im���-Fx��3y�M�֧�˓#��̀��I~���fA�L����% �"p��oR��fA�L���*V��4�04�jf�)���wC���>Ft|��q$����Ib3o#K�;�=M����hJ?���P��I,q��Y���	v���]�%3������0|BHq�_AF�6��9��ܰ�Hq�Ӯ>.��s��t]�%3������0|BH6A��fmO¶��r�``q��:{��� <&�M#���}�|��p�Ƕ���Aؿ����Uh�*�bh�H�)�l�����?یC�1�9���9M��ܠn:�2O�R�<�Uh�*�bh�_��f�/\�P�����\����"t���}'�v��w��SP}�E���[�#&�aY�eW/Sh��Fe,�)�ǮH��������ū|rI��zm���e���ş�z<�7'�x���|���s�����U밌ٓt��nG�X��%z���!��Tӧ~z,2�wÚU�	vn���D��/-�!ͪڕ6 �3RmRK��A/;���FH/Q����؉,�L��m>��RN#c�@�4��V� |���nNz�x�J�IZs��ZpK2��G'��h�x#�L_�(D{ͬ�y����"��y&�`%2
0m n2ϒ�ȗ�tVFɑܴ�G|�gL,89�;xI|$���"�|�E�`A���ٿ�,ܪ��G���W)�K��N����l%��`O~�thq�G��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������R"���c��o�$�a�Wц�>�1 T�V	�tL��	f�g���Z��	���
�Ɗ��W}g�!�`�(i3��k��my��xǀ�l%��`O~�thq�G��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc$��+�{c"G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F~�?|�[_wȵ�e�kY��Y+]��=W�֯�^��N�&��)��m��[4�l3�7DY��SV��8Q~/��ʓ|�e���O�q�Y�N %c�G͌4s+�nyYB�Aiy�!�`�(i3JHn��z�������'��%�a�9���Ő!�`�(i3�b9������ճY(1�*_��h��U]��!�`�(i3l0��F��j���^B_��+kG��!���Ёy!�`�(i3%Ah�%4
>��XP���O�w2p��AJy��$]\� ���3�ҺIÙ=�Hm�ܾ&
/=3\H�_N��-Ɇ�Q�^�y�zL͊�q��p�ΆsxI��'�����k�r�E����F�'n�^0o��vK>��5����`KB����4�"�,�>E����\�vŰ/&����͌4s+�nysE;f�Q�!�`�(i3JHn��z�����)���%�a����KG(�!�`�(i3�b9���mj��mi�d1�*_��h�Dӿ�N�!�`�(i3l0��F��jT�����N(ba�7���J��xi�!�`�(i3%Ah�%4
>��XP���o�ؔ�W����JBfϭp� ���S ���3�ҺIÙ=�H޷�LsP�=����Vʭp� ���S�Q�^�y�zL͊�q��}�-�w���I��'���gk��E����F�'n�^0o6��U�x���5����`K"��+&V>�"�,�>E����\�v�����/٨͌4s+�nyIPDa��"�M��JHn��z�_c)���8�o��Q$�"x���$�I��'�<;e�����h����]H�'n�^0o@�~T�@��5����`K�%������m�&1�]�!��	Ǹ�y85��L�?Y*�z�WC��"X��[�|���M�n3�M��?T��n	|�5����`K�%�����KԈ!
7�]�!��	Ǹ�y85��L�?Y*�z�WC��"X��[�|���M�n3�M�������k�5����`K����Ct\�|�f�.J�]�!��	Ǹ�y85��L�?Y*�z�WC��"X��[�|���M�n3�M���Fh-U��;xI|$��n�h޶��	�̵<x�iJ[�FUԥ%���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�ħƿ�9c�1��8�h����,����^�V�.�	g�y�gߠ� �`g���yퟻlA��4�	g�y�gߠ� �`g��q>?�=+��r�1�L�Xڈ*-È���*+��r�1�OG�mA�T��2���-*+�m2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�� �W9���+��l��b�"�݀`A�����xM�� �bRw�����IL�+���+n��ڃ<�8]��C$]b�<�@]fJ1���#oVhd���=�^~_|����E����F�+�/��f����U���޸�"]�IM���E�>�VT��V�&��'u�Nh���J�|(�����b���=֑�	KU�kMgKWJ�ɕ�h�4���N�����{�����Mi�$��>Z����NIi��N���o��thq�G��2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR@�/-��E���1�/���yퟻ�xʸ�f�����oP��S���Hhqu!���5�Nn���4L"�+�va��2{a�t P��;06F���b�<o�nïi�q{�f��a��4�6�t��;06Fa�T��r�m��U}�	�~v�6�(UzL͊�q���Y�egN��t���6��^hq��:�}0�st&���\�vūx`��:���Ϥk�;��|B}ø��y�w8#�RC�G�G~��6�A�7�s̕O��S�7�я�e�=��E����F���8�TP!�`�(i3v��K.Ū�C���D�rcJ]�0�!�`�(i3!�`�(i3�b9�����9B7��Qއ��0��]��cg�ų��'�oD�!�`�(i3�Q�^�y�����9�!�`�(i3�	O�\29����:V����	���]���/�b
Dy�F��m1G:D�;޲�R����fF x>H�|�!�+�"�,�>E����\�v�!�`�(i3���(�����Z8"�|o	���=l!�`�(i3��Q]� _�rs�i���H��	/�q3Oe}��&R�H�!�`�(i3�n`5�fK��0z�cUL�ڿ�|3$uJ�ܭ�PǨ�o*� 7�v�ԯ����fbK7͍��|��W&":��!Ē���x]��n���B>X��
 ���3�ҺMC�^�.�]"�,�>E���e�� �a1�z�!�ݢ�u!��+_�i������04Tq�`�����L�+P�X�;Qn�Ix���!B؀^N�ڵ5�Gi�gݚZ��a!%Ah�%4
>��f���T,�;C@�������E���7D�EIdQ�;{�rҴ�i+'��\�v�!�`�(i3y�Er�)=�ᏅN~zʎ��gB?/i�M���%Ah�%4
>��f���T,�;C@�����S-���r�a�n��W�ɝ��c�D���a��!q�N�g�]W�W����p�N����S�*H���	��<��ݒ:�NMe.��nrm؊(�-9[c9&g2��\�b�b��J�<��F�w�]��Y/�?�^�d��d}7Ê7�E�4'���Xw���\{�Sծ��[�$�o��C!T*�q���U�̬���	p��Z�-�챓=/NN; <��HT� s�yze�Zv�o��C!T*�q���U�E�KZ �7Ŭ�(�a�肢�{l�f|�-�`��8�4�%��mz%���=a\ո�k�K��l;U�2y�������5	��]�!��k��v�Kp��}�G�@����1�DX9dcY_}�n1��{l�f|�-�`��8�4�%��mz%���=a\ո�k�K��lLc�Ո�D2�����5	��]�!��k��v�Kp��}�G�@���r���֠�k+�L�)�{��{l�f|�-�`��8�4�%��mz%���=a\�&'UR�q������3���R�����+xk^�����0It�Yl���#�]�!����KR�3�[i�`#�Ք=�� Ɲ�Y^�i(�K�����b@T�!ϼ�Ávƥ4�,�:�'t��t�W�lT[�HF x>H�|�Wǖg3ȓ8���/�A���0v7�^�j����o��C!T*Y�{'%sAX���	qu�=wx4���܂A���0v7����9hv��o��C!T*Y�{'%sAX���	qu�=wx4���܂/���:;aR[�T�.�W���1��~�yD݃e>���K������j�RiP���uV�f�YcW	�TD��ό���.�RiP���uV"��J���TD��ό���.ӵ�8�,wO��oV'$��TD��ό���.�	'���~Q�<���"�s��Yȑ�n���H&���,�v�?Cc0�욁�o_��ü~���U��g��U-�e%��.�u��.�#U���Yl���#�]�!��	Ǹ�y85�΍y� I�M9)�����m"�7�����ʲ1���"B��$I��w��,����Ȥ0���a�D�"B��$I��w��,����Ȥ���_��"B��$I��w��,��xc�l��m
��5�(�����:x�V?W^�d��d}�����
L'���Xw/���:;aR[�T�.�W���1�I�$�}�[���;�q�#7G#+������z����A�b�*܋���}7���x�|���*Yl���#�]�!��k��v�Kp��}�G�@����uO����(�=���j�9��(�
t�ژq���U�$��	�fѥ�[���В����m8�{-\��]��C�yG7��6�X���Je>���K������j��J���۞h�G���d�;[��TD��ό���.��J���۞h�G�R�����u�TD��ό���.��J���۞h�G��G�¨z�TD��ό���.��J���۞h�G�Xx�Hu(�TD��ό���.��J���۞h�G�x^��+�v�TD��ό���.��J���۞h�G��!\��X��TD��ό���.��J���۞h�G�t�Ja��TD��ό���.��J���۞h�G�W�4�2�8�TD��ό���.��J���۞h�G�"x!P�Z�TD��ό���.��J���۞h�G�rv�Bj���TD��ό���.��J���۞h�G�X�fF_>��TD��ό���.��J���۞h�G�0���B�t��TD��ό���.��J���۞h�G�u��gB�<�TD��ό���.��J���۞h�G�����<w�TD��ό���.��J���۞h�G�@�yz��TD��ό���.��J���۞h�G���\ͣrQ�TD��ό���.��\�|b�����R�à��(�
t��Y�{'%s����j��0Y01�������V�O
�_�Z)������
j��qZ1�!�#c<��z��}�0z�cUL<�s�g�?�Y��Ș�Ze0G���a(􆿳��!���
faՊJ�,�w�<~t�yHJJ�5q�P ڨ��S���Q�V�ɶ�w����yퟻ�xʸ�fH(Ť"Of�8#�RC�GAPL�hN��5����`K�y �谝��X�e����yM��$��XP����+t���P�����О.�8z����&��$�RmHX���i�k�Zׇ	JHn��z��k"����_<mDrW�B���BC?T��o+W𩡛�5����`Kˊ�jJ#�}�����О.�٤\��X���XP���e����!�?2^�9�o+W𩡛0aD*������qq�S���G�M���5����`KhS���ݛ����f�u�|7ʽ�'n�^0o�q�O��I��'��3k1x��Tl\�m*�Q�^�y�zL͊�q�����"OZ���b\�#��ucZ{� }�Ri.����l�����N���!�`�(i3��Q]� _�rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'0i���crp�w�Ve�U�ԝ5�͌4s+�nys�;�srs8y5��D<��$e��]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s�ui�铤8� �w� G�"�|� }�Ri.����l���X�=1�����
�^��j"��Q]� _�rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'�k�/��O�w�Ve�U�ԝ5�͌4s+�ny����,jG�7D�EI����I�O�]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s�g��K�n��8� �w� G�"�|� }�Ri.����l����S�*�O���Y�
��Q]� _�rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'�����DM��w�Ve�U�ԝ5�͌4s+�nyx�L|����-�X���o"�,�>E���]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��rs�(�̴Y�{'%s/^)i�cϤ8� �w� G�"�|� }�Ri.����l���XB��$l��P��N��x�o^�Y�rs�i�H���N���w�Ve��t_-Z��T�\ ��QD� ��-a�vݝh�c�A�L'xM�0�5;�w�Ve�U�ԝ5�͌4s+�ny�y��P�p�V��O"�,�>E���]�!��	Ǹ�y85�|읯2�9�G�"�|��ߪ��wZ�n��[��{_8�Y���˂lq��r'��i�B�J@�l�s[�5����`K��D�	a���Ӯw!\�8䮨��ekW���I|JHn��z��ea���4p���eqd���w&�r��VYW\�����[!�`�(i3%Ah�%4
>��XP����~��84Z�Ћ�l�TE�խ������S�0ů�x� ���rs�i�Vw�C�-��0#�tC%Q,!�;��
r7��(*h�Qf�kCH`=Th=mP��T�͌4s+�ny\D}��^��ٙ�D�s^E��S�Z鎬�������(���E�̱!\Z>�
6������+$��g��U-�e�v�W�G�[�^�������-the ���mh.�]����GC.�|���~��H��efm�0z�cUL���a��<mDrW�B��"���PB[<b�P�`<����B��٥P5���rs�i�H���N��C�X<� ���B��8�R�Z_.΄x�g��	��S8��UV��\Ƴ�r��Gh�Qf�\l{�"7�sa�vݝh�c�A�L'�1�d��{�ʬ�缆�YW)��͌4s+�ny �Ǧ�_@f���_t��R��XP���x���: �&�(E�{�ʬ�缆P �8�-�U���L��$�y︁��ڨh�ϣ����l����S�*�O��a.��%h����]H�'n�^0oP�M�'?�S�5��'!(��`�\s�I��'�D�ԗ�CW	�h�b9���O���2�N1�*_��h+�I��|E����]�7��Q�^�y�zL͊�q���ǹ��L�I��'�J���̯u)!�`�(i3�b9������ϸ�t�O�&����4a�5>.}V�� -����]�!��	Ǹ�y85��L�?Y*�z�WC��"X��[�|���M�����Ct�O�z��l =�������A��J�E���V'/7s�9���o��S8��%�CF�I��r��Ȯ��ߊ��H�R�?4���-�ܪ>�����K�Q�f�;�>)ʁ���f��Y�{'%sgeߪ�{ ^�x~�(vi�t�c,�q�T�\ ��퍥6� �iE��_�/`C�|�dz���$Z鎬����Z��C�Ջ�+vTń7���*��P�Y�
�d�٣�����6>��w"�_y�=�ꖯ�y.��&��ࠅ�ﻋ-�����S8������ۓ8���/���J���_?��]���g�(�[�*!�`�(i3��Q]� _�rs�i�;���fwa�\h5&����8���/�l|�*"k���(ӈ��h��P��u�һY~����I���a!�`�(i3���+�J��p�VU��J��'�����1 Ҏ�������Z<:9�-{$�����v�}��Iћ<���E����FZ鎬�������(�����dH�L�p��HM�e��Cҷ��e��'�����1 Ҏ��7_]�4"m�S�K�Q�]qE�&��R��һY~���L.bC��!�`�(i3���+�J��Y�{'%sAX���	qOƋ.]$�t_-Z��T�\ ��w�vܖ��X5�:��o� F x>H�|�Wǖg3ȓ8���/�-�',��|$]�6�����_��u��th�_ME�v+�	k����tp�p}��qΎY�'.������մ�g� �P��}�/Üy�a
�i�uŕ���&�&�IE��K�L"eOx���'RFtI��&� }iIB?�d�٣��c�A�L'!_���#��t_-Z��T�\ ��w�vܖ��X5�:��o� �w�Ve�!8���\/Üy�a
���"X��[�bwKL�G�"�|��5��ݦ,qqݥT�Jɇ����$�x�Wt��Q]� _�rs�i�H���N���w�Ve��t_-Z��T�\ ��w�vܖ��X5�:��o� �w�Ve��t_-Z��T�\ �͙��D������ΰa1���5�'.�!�`�(i3�n`5�fK����3E�Y1f����٭(��K=J��(�n5j�?�T����g��n`5�fK��0z�cULCx&Z�����8���/�l|�*"k���(ӈ��h��P��u���v:,{��`\5
��0�%ً��d�٣����>2�p�n5j�?�T�^'��s_ㆂ`Z"�A�?3d�!TZ���|�E���I�u��ʝ�Qer;y��^u'�wp]Yy>@��$n�m�;;���գ'���Xw}a�֧a�A�zB��݋����f����{�&\��n(n)6�0�4��l�7���H>����斣�������6p�k&}ǝ^3�n`5�fK����3E����}7����a*`�(o&��͎�e!�`�(i37L��1�6`�v_�w\(��gz��}�9���P��r��c�@#$Kb�i�)6yҌ��7s�9���oC�M��N�ې�7j�5繁�~?R����I�
�2�� Ϳ�$�<ͧ�:|�*�za�Hj��7j�5祐 p�;H2��I�
�2�� Ϳ�$�<ͧ�:|�*�za�Hj�(�Y�MMoߙ�(ml���d������ Ϳ�$��0z�cUL�{���7���ԓ�a(􆿳�����0omwj���dDq)�{� �""�,�>E���]�!���1����m^��PN5|�B"��D�a��zr,/'���Xw�����C�pzl��a�G_����\ό�������n`5�fK�<ͧ�:|�*�za�HjWT� �`�o$�x�Wt"�,�>E���]�!���\B��Vm5��i�����`�����+�����+�J��p�VU��Jm�QA�Q* x� Y���틅&�i2]�5�x���1R�W+`�x�oP��@t��4�u>�[�9q�Y�{'%s2�ew���o_��ü~���U��g��U-�e5��e6²���R�:���g�!�`�(i3��'sT:vSk,��-�
��LQ..�e+X�&3]�&�F�K7͍��wAA�Ɓ=<�W�.�P�(o&WQ5�xY[�uB�|���yG~F���g�Ww�[h�q��!���\���Ȑ�'t��t�W�؏ 4�+�{_8�Y��M��)=໺(ӈ���x|}�|0�D6}�������2�k��in*�k�����\F�^�	E��߅�'e���婣	���U�dN�<@Iv�H�_��Q��b�z'hۉ)�5�c*�{��K�Q�J2)V!�`�(i3!�`�(i37s�9���oC�M��N��y4:��P�΁�a�n��!�`�(i3"�,�>E���]�!���1����m���I�@�!�`�(i3!�`�(i3зq8�Ј'���Xwa'�<� \��͡��!�`�(i3!�`�(i3��Q]� _ό���.�pzl��a��X�~׫�焃:p���6��N@u�Y�{'%shM���V��>>�%�/��ㅬ���:F�X?�g��U-�e�_|�<�Ԯ2X����t p� k��*4?���]�!��	Ǹ�y85��A�'�/#y�,����	�H�ɂ��:F�X?�g��U-�e5��e6²��J����$�䯯M������/�C��c���d�٣��c�A�L'c�y�l�jO�DW�IP��N��xL�ba���"X��[�z�C����G:��7��3���Z�k�X�zBg}1ʾ�!����� Ϳ�$��0z�cUL�ڿ�|�CL#�fڸ����@�ս��'v�aW�Ȯ��ߊ�R�wX�՝�E���8�Z:���6�D�J�4'���Xw�j�7���.��y7�N��b��%�����+�b_Ma�~�Ǔ8���/�p�.K5B��R���,.��.��y7�N��b��%�����+�b_Ma�~�Ǔ8���/�a'�<� \�&on��l);�OA�uWSx�lޞ��rs�i��-�ѧs��ʟ0B�@C	���{;-;*�7���Ȯ��ߊ�R�wX����츕�)��d�[�+�dJ�ܻ���������e�1��.);X��Vo���4�"'ɪ�#́�V�,I�Q�,#a>l��Y����|�=��d%�Z9`h�-����M��$4N n2ϒ�ȗ�tVFɑ�k���8�āGN�~_�/����i���w�6�����́��vn�y<�f��`-�B�l�2��%\EΎ�t%>^��?�y��hL5ӥ����c^����
<ڑN���2�A��1��R�9*�eaA�|j?�d���&���>E��*�(��z�¿-ǂ,yߊ��b,�a������)�}�����T��.��W����t�.�!�8�}�\���;A<�SNp>�3������"h���ƅ5����5�`��N�W'�o����f7����e��x����#E`D���$G�	P��?[@S�CZ�~۵�q�#�p�	;�0�e�n�xdɨu �䆡X�dr�jf'��H������V���
���F:_ʣX`��_/��IC:GMG�2�3�A�E'����>E��*	Z�~(jm�7jl�N�Ar�/=�N�}���X	j�w~jiǎ[��S��_�:�R��h�4�b"����gE���Y(��	Q��H/!�Sy�+�z�}�-�%Q�a�4f�+�Z�{�b7�-�4T����	��,��<����r�k�,��~��U?'�����ٴ��{�G��ͫ������:[ۚܖ��`�[�	2�GF�&���#VW�GaAO'��7wT�,���P�&`bH$��>��L��$�I��i�j~>�Q.Ss�@�������-R�X��%�VB�=����R��(7�
��o��N⃟g��|"u8��d�w(�`��l4���/A� e8�~���db�_��n����L��tVFɑ�����n2 e8�~��-d�L����i���w�6������<�䛄�� e8�~����gľ�W���dx�b�W(��	!nR�*H�a���λXθ�����Ƃp��Sr��n�"�rNy$;=�@俷�v�������\��&z�0��E�5�JF)c���'7�*|��G��U��t�uY������p��V�(�\�v��
mGԧ
s���7���=�V��E�&����f��jv�!d*�[��&�[}�1���V���~�L�{�g:������(5;|)f��X+��f�������~T����H&���'��N��i��\#+��S�V�W|�B�I:׷�Fi�k�Zׇ	JHn��z��r9�3��*���3m��U}�	w�v�����zL͊�q���19TH��@���U@���:��F�j{n�}�R �i7�sp>���=��s*c�r�w��*�T�P!�`�(i3��{l�f|�ό���.��g�rz[t�E����F�ҋX����@�ڗe'e'��ǩ������I��w��,c�A�L'̙ch� 5A�
c�[���ߪ��wt��I`��8qTmI(xe�0
A���g�Lc!M�� ��P�l�U�,/����v^�n����o�bz@�o	�Au��b����`m��';��?2^�9Ͱ���*U�'n�^0o����y�]�{G�3��!�`�(i3%Ah�%4
>��XP��ȯ3k1x��T'��$������)2tm�c�oL�`:��Q1l0��F��j�mV��5f���=��s*c�r�w��b��	��碢FҼ�^I�ҋX������S8�l��`�p��HM�e��`y�����˪XkY%T��BPS�)37J*u)T{6T'`�<E�dh�o��C!T*�q���U��3|�&��J� dC
kS�)37J*u)T{6T'�
���t��o��C!T*�q���U����j��Y%T��BPS�)37J*u)T{6T's�yze�Zv�o��C!T*�q���U���~JFNǑ����E��@IE�U��w�B[��lQ�$�k\_x���� �~��Z2��l
OE�<�x��3����Hhqu!���5�Nn���4L"�#W��xW�Kg!�h�����7�$�G�j/����X�e��}c���G��m\Ӓ�qܛ�	���:�UU�39M��0�d�Sd��_�a���n�|W x�Pw��d�(ߏ�"�nT��z��uWU4y5=>F/ġ"���Չ-RW!�՗"$p\�>���S�w҄�^��(I�>'����	4T���\�nƨP�ʱ:��Ԩ�\�"ߗtl%�]Y�%���Ádo�d�x��u�5�h�br���lpda���?̕U�/j�g4A���{0Yafk��r.y����nL���~C�V�T��a׈Eg#f�z�q���<�{�!���"�ֱ��R8v��j.Z��$�sӢ�]3�����c��(r"�o�Q�E���dZ�雇�p� o�v[�(!�lV�����9��S$�xx>���nj�&3H2+lH*#$��}��r�7l���qs=j)�0�� t�!���Wn�d���T�OÈ��{3{a�T��r�m��U}�	�_ק_��e���R?�6��'�|,kW�A��ˮ��V�rsSRątG��2��ȫI��2��e��a�8���m�M��nO���$73���'���)�4�GAs`�D�dl~�)	D���$�,n���A���c\����(�a��;�<�� ���2�jE?dSծ��[�$	^����ξY'#4��e�ά@�ș�I����~u�m5��ޥ�}�gazy	s8R.@��H��~Ů��D!����ހ��g�R�N�ގ�MX@;��I�H��?5ǺW���<�K�kσ�a��R�4�}��hw��C���"BC�I�1X����w�d ������R��Q�C��1Քb�<2��]��I��o=�<*��
�]v���!�o�fy`,��8����^FG��a�v����Z<L���p|j
��s�|���죆�����w܁ZUz�@E+��nw��m�x�Z8p�nrm؊(�y�uD#�#�!<��f���f�;�>)�:_~�0�-�캧xӍ.������J�F+KK� ^���PG{��_���wE���B]DWl$�`�]
���bψ8<�!W���2��h"r�����NFsU۞h�G����T���R�<lͬ۞h�G��" Y� \���I�&�`Wq�`AS?�C<xWY�K��e�Igg�R�@�3�0�DZܤ�jM��3�}�v��	'����'�SS���L-�yC³�h7�a��c�,�[`�B�!�e�Զ��,�qm�c�,�[`�~$��q�r/�;�H���o�O.���	�i��#�f�;�>)�k`�+Y�r�캧xӍ.��,����«��	'����'�SS���Z\�i�æ`NR���c�,�[`���K��+�rF)���X�3c/��!LH��3�f�;�>)�Q��S����	�i��#�f�;�>)�Ĉ��^A캧xӍ.��k�jZ"+KK� ^���PG{��_���\��K��]DWl$�`�]
���b��278Jb���2�����ǈݻW�)�۞h�G�>��grc���R�<lͬ۞h�G����r䮥���I�&�`�̖�K �?�C<xWY�K��e�Igg �%���k_�DZܤ�j�]��	HeIYv�(�@���2����I�}j�Ez	*HD{۞h�G��������a}�%h�/�<���Z���p�VU��J�-N�W�Z���Y�{'%s��s�X�O��ςy�н/v�IX0F�M\hꑣ��P��Hǲ(-F��� ��b�FP&\�R�&�-��LZ�|�b,�n`5�fK��0z�cUL� ���Q$]�6���p��HM�e��`y�������v���д,1.��o�܁#k$�H+e�{'���Xw�j�7����o_��ü~���U��g��U-�eJҪ��D �k]��Ĳ�;R���ȥ*�sk��<�
�dW���ֈ��tX��Ӧ�Q=�=y w�⽒�PUaB�s�{[���G���ӒJW�>�ܖ�4��x��h��B'� �����T�غ�Z��s��u�FR�Gp&��fF�5.]����U4�i�x��h��B�f�6l�}C���a[SM���5��F�ύ��mCt�w#��@�O�!���͔�a6gB��{�=2|�l<�K�旼��7X��^w�̀	'��h��n���=
����l������|�Q~�4n�Q2�������C 1]qE�&�.}�I�̆�U�J�J��JT_���y{Kg��C���a[S.��o�܁#��ޞ�~*Ż�&ǥ�̻����.�fF�5.]���k_���b_!2�͞nOY�N�zS�(�xJ�|�S�	�j�����Q\�_qB6$&�������Q3��Bd�Y�k���;��-�F^�M~Ɛ"ǩ>�)E���Z�� ���K%��e�=�#�vG"J�CJ+T ?�7r���g����,	S;&�+K���n��M�60��g�0�uKK0�RS�]
���b,IE#N8��ð��T���YIt�K�~V��=�[<�����M��X��At���3�l��d��JXl'�&�P�2�PUг�|<�D�$0��;�H���o4Go�HHm��1��X��WG ���K�"A���.���G?���{Gyn��@�a��W2�X�Nb�J��B��O
�_�Z)����ג�rw�&�z<aSm�6��`4�04�jf��ܐ�}�S��/:+�e6j�"Hs����i�A8���9�D���g�b�^��\+��%S��P��}+80�o�]��y�߀�����Z���<�a�sN$ug�W;��|B����_0���"�u1Tb ���+���Ã�E؀��<]c�,�[`��ᾮ$�YZ���������K�۞h�G���7?7��I/��\];+�ܴW�~p�ܩv�iIM�j���\�����h�Z��	�IW}�y���,�1ʾ�!����o#�o�l_���%}��s��U;4���^a����HŹn�軑��r���/�ciJ�:��er?G����Oam�i��ċ�!-M�O��~��B<�q��L.bC��U�gQMf�Ʀ�|þM�I�=X�����r��Ȯ��ߊ�u*w�A�X�H�u�q0O�*2t�ch��KV� �Ĥa�	�+4D@�p�U>�tf���!���ڽh���[���8D#���i@`:v�eQ۞h�G��#@�h�R*E���&�Ut�\�� +�,��T^���^%�VZ�$~p�ܩv�ng��	T��5ߧE4��rw�&�z<a��N� φ��<�6��V�4��5a�/`C�|���K#i�Ʀ�|þM�`�1v�-�/@[�_zβr�v������Y�hg�N��Z�H�9 ���
�8��рa��N��*3M���*%C?*����l[j6�z���D���0�j�J�Ñ�����������g�R�"Ì�s��X�e�P�����`�B�I:׷�Fy�XZ@po��*���3m��U}�	��,�{�'�3�$ �#^�Vn���v_�"c�PƐt
�20)�_����*��Y~��`�J)����9	�(f���5�r*Iީ�4+�A!��X;p`�Z�^6Sծ��[�$���d~lr��[J�c�,�[`�u��s���6�ς�(�D�0�?����N���a\�î�����Q\�_qB6$&�������Q3��Bd�Y�k���;��-�F^�M~�pgL���_�?�d���&��l����F8�iE��1Tb ���+���Ã�E؀��<]c�,�[`�{��(:/�b�&�q����}�b�����J�Fbݙ��N�g�c�`�%��ɰ�����*�݄���K7͍��|��W&":t���3�l��d��JXl'�&�P�2�PUг�|<�D�$0��;�H���opwI0����1��X��WG ��F�����8�iE����8?"��!�;����OvEZ��U�&�(5�;2�f�;�>)�ӔuP��N([��}qn
V~$���d]m�B�/������T�b���'BŉB������*Tz%�vѽ����Uh1ݵp�!���׏�����MJ�1���۪	�}a4�����l����F8�iE���x2�:����ء5�訖�#H���$�MN[;��|B�K���&�Cߋp{T��c���,�\��{ElCg?	��ofob0�۞h�G���w��z�=k�Rm���8Ơ4�ܩ"۞h�G���7?7��R*E���&�j!�\B>�jK�o[���[�2ټ�mˊ��ձΐ9xWW)��~?R����I�
�2���L����\9�oA�d��JXl'�&�P�2�PUг�|<�ɐ�>8�co�v[�(!쥭*����	D~��n�&�;|>r:w�:��er?G��7Wx� Pabݙ��N�g�c�`�ɐ�>8�c�"�rZ��.�uO|&�9�r�I�;3�p
��a.��,	�g��WN������)<�-w�|��qĵ=)�7��B6Ji����|���!9�j�m�����N��4M̍����5Ɇܾ�]��	He)O,�rە�f�;�>)�-m>c.��{t�Z��P��3�Q#� :a�	�+4D@��/�ciJ���z 7	B>�b��O����~y�
3��0�ǳ�ȕ<dh�}3d�jK�o[���[�2�֚���,��Hp9��Ԍ��Ǐ�c���w�I�7ݟ=�NM���ɛ�?ө�&�(5�;2�@�a�����be�vҜ��)P�N�g�c�`DE8k �Υ4^��)�d+�����q9+t�}f��1�x���~?R����I�
�2��f��U/��.�[ ٓ��r_��mԌ��Ǐ�c����3�6oݟ=�NM���ɛ�?ө����h`�CgD�|�݄����Mv!���xx(�i��/RŻ�&ǥ��a���F�LFC7�5$�)�vx/�k
�SR��Y0R�ne�>�H�ܕ6��HHD�u���&.)+�ޅn���(��h�*蓱Wxi��o�bB�۹�D����=��Y��RJWz���
9�5ARL��׿"aj$�b�w}P�
���(�����d��R�Q��=�ƆR�(o�Y�f���'v�qB���jK�o[���[�2�gu�}���<�f�;�>)�-��a�A�so��%���;�N�cP��&��h����E�F6���Wz�o�3p�60���!��2��J�J����3%E��_��=��}xsEqFM���K����x�l��15�r*Iީ�U����W�!�`�(i3��a����9��>�������q�}hfQ���f�d&(C�#�7#^�Vn�zy���l�?2^�99h���<��p&Zc��g}Ю�0$�W���AO��ē�����1����S�0�b��Q[�f�8T��=���� �h�
Xק|"��\Vڜc�,�[`�Z*ik0��0=�!�hj�|"��\Vڜc�,�[`�,��΋�ߏ�sH�
9�d�(�?��~?R����I�
�2�#/P��tZ�H��S����QM@%�
6u��'Kl�����.;�<.�2� rѻ��S�L(�y�}��;����<W�X�ﵤ�'D�<������>��}��lj��
�j����H�A���������KX��ik��dc�@z�ׅ�ؘ�X��WG ����[m���~/�9�(���[C�/������j@fq��]^] c�j*�/i�D�]
���bۖܧ�k�%����}7����a*`�(oV���B\�R*E���&�Ut�\�g��j�n��뾦��"L?���)@�-�� ݟ=�NM���\n0�8�׏�����Mx(�i��/R�������a�U�ے
��]3;�Lmv�)5�/��-0��߷�ˎS�W���tkU�#���.�����?�#�6�f���!Qr�g?	��o`
��3�l�g�0�u���^a����HŹn�軑��r��4M̍����Y"�g�YZ6��HHD�u��'J��l�o=��i֌]��	He$(�2�ft+�f�;�>)�;��e~]1bt�Z��P��3�Q#� :a�	�+4D@�z�+��pQx�(^i��֚���,�%][��"����@�{V"s�ֵ�݄����Mv!���x�5ߧE4��J�1���k_���b_!2�͞nOYN
,k��"�Z2k�VKY�_%Dό��סزN.�Xkez��Ck�8'��d+�����o�½X5�g�0�u3L�6(��dM�+���T�>���({")8�*IO��(����׹��˸$��C�r��T!�z�د��̓С�*�WE��by��Y"�g�YZ6��HHD�u"�T�B�Z��4��)��P�>�n5j�?�T�P�� Rܡ��d���<h)�!,�!���^a����HŹn�軑��r��4M̍���?��ㅍ7b;����R*E���&�Ut�\��,2�C�����d���Ą�Ĺ�,7�cL���	Ǹ�y85��֟��D�D���P�ħN�g�c�`�9�d�L��s"�k
�5��)�rbJ6�~��Jtat�r���N�g�c�`����m��:��A��+���4L"�ɲo�I�xg�~p!ۓt��p�O%�70��G�F���"���e��d��Nt7��?��w|{�ۚ�7���.L��h�T�W��S�� ��9�Q�#�ͫa���n�e�[7�w�sB�ƛ��pP�����d�n5j�?�T�P�� Rܡ��d���<h��Hp9���5ߧE4�훬�pP���Ǻ6�(c#�ͫa���I˒��M �ҋ�;K���L���4�04�jfx(�i��/Rh�x#�L_�(D{ͬ�y�4����W��IW�oQ���`�A}�/6�o8:4�;8I ��*��]��s�6e���im楰�z*��['D�C�k�a�	�+4D@S���O��zB��݋���>?���{��G�����
�]W0�e 6A��c/�w#�ͫa���n�e�[7
$B�>���I����~u%J�bb��|k+Q�h'�Ȝxڣ9�$���>��o��%�C�5��#���+�9-�i"'���Xw�j�7��FZ����^��h���LX��WG ��2�t�N��y�R�QY`�CgD�|���$�!$Y���@�}%@�`�4��h�3��'c�,�[`�t�)
W�k��
�!���i��ċ�!-M�O��~��D�$0����=�����Lj1���7Gvz8�uX��WG ��Ĕ�.p�1��zB��݋���>?���{��G�����
�]W0�e ��Hp9���q�;������\�2���.Z��'!�`�(i3�kȹj F~��h�T�JDn ��a�'���*�e��@���=�����Lj1���7GR�0�;"��9�{�n�[O��nD�%�z�J���o{��:�N�#�@j��{�`��ҜcZ�����=�<�^�c*o��ܔq_�pk����2%g����<-����R��n5j�?�T�LW�_��%3�o�:�>je`��@d�,2�C���l�yi��L.bC���Ӥ�bϩs8y5���PV�q�-n
V~$7���.L��h�T�D�ԗ�CW	�h �ҋ�;#P�j2E�?�o{��:���m4��0���f��J�a$�Y �=�<�^�X�H]��9��6�j��n	Y'F�0V����x���g��̙(�j���%�z�J���o{��:�N�#�@j��{�`��ҜcZ�����c�Z�~�c*o��ܔq_�pk����2%g����<-��ic)�̩��ɛ�?ө�e��@���=�����Lj1���7Ggx/Ҁ{�-M�O��~��c*o��ܔq_�pk��=��hX��9�{���J�sׯ�ɛ�?өW�{OEׁ��q�2��Kk:)���2��D+���4Y U�����p�zB��݋����f�� !# D��B�R���>_�c*o��ܔq_�pk��=��hX��9�{���J�sׯ�ɛ�?өW�{OEׁ��q�2��Kk:)���2��D+���4Y�q9+t�}�P�HS|�4�04�jfJ�1����s��U;4���r}�L��Ώ<�?4Ck�8'��d+����}�{LFv(�c�,�[`��� U󤹼�j=/x9��c+
�i�l-�	�yH@�
@����=7�}|��	��a-6�DaH(Ť"Of��D7��\�b5;4�<Z�g
aC��en���o{��:�N�#�@j��{�`��ҜcZ������\b��z\�Q��TXP�e�g�6�<+sӑ�fg��n5j�?�T�^'��s_ㆂ`Z"�A(sB.��Hf;[���7���.L��h�T�JDn ��aP�d�����a��R��q_�pk����2%g�p�X<m��J�1����ݾ-/�uu��ڿ׏�����M��ܐ�}��t�l��뢂�ʆ&oA�\ֆ��p*��2')�F	K`���$va@)�	��x�{�*~��Ez���rJ[����0+C�t���� ����!J�/� �1x�it��l^�28�v����l��H��efm�0z�cUL���ޤ�Y581���5�o�N�g�c�`��QU�+J"�=�<�^T۳�͕��(̠F���%J�bb��|׏�����M��ܐ�}��t�l���sȸ�"rR!�`�(i3On�������Fz�!�`�(i3���w�Eo��]�U��!�`�(i3oW�����Ƹ.��v�!�`�(i3}S����inca߫r!�`�(i3�&e(r�
=�4�!2d!�`�(i3�1'�b���l*�����l*�����l*�����l*�����l*�����7���Y�����Fz���>�&?(�1�f!�`�(i3H2���b��(�[�*!�`�(i3!�`�(i3?��h�|�!�`�(i3!�`�(i3&�{��x�l*�����l*�����l*�����l*�����$����!��Ƹ.��v�!�`�(i3�n3z(!�`�(i3�ng�[�^!�`�(i3!�`�(i3!�`�(i3?��5��!�`�(i3!�`�(i3�R�
D~��.���{	RK2�����Vc2�����Vc2�����Vc����:��Ƹ.��v�!�`�(i3��_�/?���d����Ѕ�WX�����s����t�q��!�`�(i3?��5��!�`�(i3!�`�(i3�R�
D~��.���{	RK2�����Vc2�����Vc2�����Vc����:��Ƹ.��v�!�`�(i3��n��`
H/Üy�a
�D+���4Y^ �7�}3�d"T��O$!�`�(i3?��5��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3Q@w�ӏ{�Ƹ.��v�!�`�(i3!�`�(i3!�`�(i3}|@�3[J��<�,U?t2�����Vc2�����Vcc��f�.E!�`�(i3!�`�(i3!�`�(i3'q�%ȗ�5��p�z8��x�?J,��j��n��&<C�3�Ƹ.��v�!�`�(i3!�`�(i3!�`�(i3�E�a��@����Q`t!�!�`�(i3!�`�(i3?��5��!�`�(i3!�`�(i3!�`�(i3_j��u��[2�����Vc�/!��v�22�����Vc����:��Ƹ.��v�!�`�(i3!�`�(i3!�`�(i3ɦCNM��FY��/�.��?��B�G�"�|��9e�O��vt�dZwIF��`\5
�1��9��>F������>?���{��G�����k��k|�5�������r���Z����Qj;b�R9�����KD�;E���D������V@Bɇ�L�C���ea�Xi��`
��e�� ��.���-M�O��~�Nv���å�12b5e��0�U+�qbp@���a�z6�F�KD�Vr[?z%CS2b-M�O��~�Ѩ�f?�R�Ԍ��Ǐ�c���w�I�7['D�C�k�a�	�+4D@�K:+>���}�b�ew�T'bݙ��N�g�c�`��L�ΪA���Ǹ��St��h�T�D�ԗ�CW	�hi��ċ�!-M�O��~���L�ΪA�%�C�5� Y!܈��u@f�u\@(H�o��΄x�g��	��S8�>���r8j�g����PTse��ͳ[�%�z�J��w�
z|�������Ʒ����V�3��yɶPі��/�Z鎬�������(����ЊҼ�<���v��H�h	OB}ә�]�Ϲ���6�|�MX����N=�rs�(�̴Y�{'%sAX���	q���x���:�M�C��Ut�\��ɺm7�{L.bC����s+N���D��N��c�7,�%����Q��������Ʒ����V�3��yɶه� �4�<rw�&�z<a��r���T۳�͕��9�d�L�� *�P�RO�?@Pf)�+�9-�i"'���Xw�j�7��FZ����^��h���LX��WG ��"��;��	=�T�f������d����1l.���7�cL���	Ǹ�y85��֟��D�D���P��K1Y�q���Ȇb�L��I�d��u��H��efm�0z�cUL� ���QVJVJ@��/Üy�a
�u������n�%�z�J��ʛ	����	x=:��\�R�&�-�t�{O�v�dfP�x;Q)j�R�c�Q��Ȇb�L�������3t���=�4�04�jfp�-a�D͢q��`�L�ʛ	���<���&�����?��zR���bʴ6 �g^�k�����aD��!C �@nk�P�U4}g&>je`��@d����b]
���b��4��.@/��r ��%�z�J��k�z��4��[�}��|���Z�^������(4ޓ���@�wDJ�����.&F�Y1f���V�@�"�<đCM��ߪy߉�m�$rw�&�z<a�4�ڈt׏�����MJ�1���۪	�}a4����@[�_zβr��S~��5��B4�����ӵZ#=D;r�R��x�K粞ƿ�Ս���:�!g�L�aB^v�Ċ֩��e��cx��Og�&LTXP�e�gh:�:g�/i�M����}������3,� �Ԉ����Ia+�3$��$#z�*,�c����Gp���������
c��m	UZ�%�!�v6��	X%+I�$�l'�7��ܓ��;�7�v�FpbO)�����Z�H�9 %�$����ۙ���-!cXp32|X�=í�����jXؤ����p�J���K��S�&T�ͪ͌<4C_�kQ����Lc�TH������7��ʒ��mY�G�В� v$���K��6�o8:4�;8I ��*�n89j��<$�g�0�uM`B�Ӑ�>�b��O�=7�}|��	�3�� �fkx8냞Ă�nF���<�W�.�P��Dbgo���k+Q�h'�Ȝxڣ9�$����3�� �fWT
Y��%r9���TLB������([��}qn
V~$8Ơ4�ܩ"۞h�G�2B�_p\_R*E���&�Ut�\��ʛ	����	x=:��\�R�&�-�t�{O�v�dNI��L'�!�ɺm7�{�I���a5C�>��Ei�a�sir�@�A��I����!G�H�E U�Z��Tx�&ޓ�TpR0��ok%O�kai@`:v�eQ۞h�G�]t����qcR*E���&�Ut�\��F�R�M�ЯҞ{��6�.2�MWgX�����vs��P�<��^NEF/H�x]o/�� �T�1 Ҏ��7_]�4"m�u*w�Ac�}���Fo|k�Lbx(�i��/RŻ�&ǥ��a���F߸��S�Ȍ��"+VqS?�d���&�ۙ���-!:+4����_pQϧp��k�����z~U�6B�Ba��;>��N� c��Yi�����>F����B�n��'���gB?/i�M���;��Qz�#g�k���6f2m�ڬ8��ٶbbD�;E��}Q'(�!��B� ��~�� ��B@XI6\�4�@���(�?<n
V~$ً���N�c�,�[`���W�XN=7�}|��	��a-6�Da�J�$����&�ߍJUv[S�d�a�vݝh�c�A�L'2Ƶ6�G4�a�T��r�m��U}�		��99j�RmHX���^uU�:�|�)�6>d�r ��a�z6����}�b�;�N�cPbݙ��N�g�c�`�c*o��܆�m]jx]��4�6�j���{Gyn��J�$����&�ߍJU��Xf��� 0��#�'Y��m�xv�O
�_�Z)����ג�rw�&�z<aSm�6��`4�04�jf��ܐ�}��L���-�/�;x��A�d�LIX�"J�CJ+T ����H�A�����'7�j�s��d��JXl'�&�P�2�PUг�|<�D�$0�y�R�QY�v��|���A�$������elk��۞h�G�2B�_p\_R*E���&�Ut�\���k�*�V1��1 ���;U"�$�|.FH�韓X�HWT
Y��%r_�1�J��]LB������#o�]�ʄ��j	5�j���g��ǻ�Ji��ċ�!-M�O��~� t��O%�x4�#�:�j�Nh2M�r!t p� k��K�(�3$uJ�ܭ��(��㽶v�I7��-5�O
�_�Z)����ג�rw�&�z<al����HZ�D�$0�y�R�QY`�CgD�|A�$������elk��۞h�G�����⚴R*E���&�Ut�\��E��b4
"Ohƪڈm�H�Nb�*Z鎬�������(���� �L�Nj������}zES���)�9�Mȳ-桞=�Q��v�灹/�Zn���㬺.Q�r:���.￺Ky�R�QY�v��|���A�$������elk��۞h�G�2B�_p\_R*E���&�Ut�\����x��,����8�e��=�u��N�g�c�`1���������8�e�݄���٥P5���rs�i��-�ѧs��ʟ0B�@C	���{[�W��g ���8D��d�Z�� bi���0��E|�,z�X
3kZ��˓#���gV�p9�5t2��� t�p��'JX_)B`����'�mH΄x�g��	��S8�4�m���=�Q��v�灹/�Zn���㬺.Q�r:��rw�&�z<a�4�ڈt;S�	Z��rw�&�z<a��N� φ��<�6��z%�ژ�(���f��3A	>[��G@b� p��n�1Tb ����IX0F�MN&�'V��g�0�u��L�4��j�Ï��	�Li4"�	��z��R��Y"�g�YZ0��3Ts"�T�B�Z�b~*��s����{?tQ���3E��٥P5���rs�i�Ǘ$� ��������-|�w�������=�����Lj1���7GXB��$l��P��N��x�4��aa�<d���u�q0O�*M��3�}�v�5�����Qa�	�+4D@vE7�MW	>[��G@b� p��n���`Xg?�=z��k�8c"<�}�e�K�����	wYMՙ�o0��{/��&�<ay�N��X	~lO+HL�hG�[Ø�;�xx�*aE�8BW�R7���so�-c�,�[`���m��J=7�}|��	��a-6�Da8�-�]/2b�e�q�]k�WM��q�݄���4m�s�I���D�cɱ/������ng��	T�x(�i��/R#k�˟ܒ�o|k�Lb�5ߧE4��\�ܢ��,	սL��$�\�|b���{g�e�?]�^��"Ohƪڈm�vdϣ�k��4(/9qy�BdQ"�&]����,�ǰH7"LTfti #�sq��N� c��Yi�����>F����B�n��'���gB?/i�M���Ŵ#����#g�k����k�*�V1��1 ���-x�<����쏩C�:k~���c~,)�z���:p��҃d��{S�G_����\�f�MX�xI@[�_zβr�v��������` �6!7:~�W��;7>;B$����D�,�H��)�u������k	D[��r������Bg��5;��Qz�#g�k��q쳚�=��20{�(m��M��X� �w���z�L�C���ea�Xi�ݮ�dc�@z�ׅ�ؘ�X��WG ��8Ơ4�ܩ"۞h�G�]t����qcR*E���&�Ut�\��=����ό�������ڙ��H�m�*,H�3w��[#M���*����	���hKˀ�P��5���Qu��˓#���X�Ȥ����A�qL2�c��mˊ��ռ+���8�׏�����MJ�1���۪	�}a4����@[�_zβr�v��������` �6!7�bh�e�,��[u+���
zz��~��"����6h�烋�ɝ��c�D���a��>I��uO[H5�N��gڟ4��&�jW� ����!Qr��zj7i�j�d��y5\����������������3��a���Cوj�~Ut�\�����b]
���b��4��.@/��r �*s���j���쏩���d�F)���+Z��\�G���:��er?G�Wq�`ASi��ċ�!-M�O��~����M騪�A�qL2�c��mˊ���@�.貣�FU�D���9�@�r#�9l$U̑�1G`3n�ea=�x��/"d�GR���쏩���d�F)f;[���J�1����ݾ-/�uu��ڿ$�)�vxe�zA��;��|BmB�ut�=7�����bw��2V�RGS��=[��uܖ��m�el[�����N�9�?_��s�֙>�5�(2�q�is��g?	��o�dEr�+��#ȕ�B�������Ѩ�f?�R�g��j�([��}qn
V~$�UӇ��ɋ� ��X�D
CvK}D�؈a������h:h_Q\�=<�6>e��0�U+�qbp@�w�&1�|���yG~FsW��/dN�<@Iv��nt=:ྵp�!���Ct�w#��@t���3�l��d��JXl'�&�P�2�PUг�|<�D�$0�y�R�QY`�CgD�|A�$����@/��r �a�<d���u�q0O�*2t�ch���5�����Qa�	�+4D@i�a�sir>G���Mg"�jw�|�L�K�p��x��_�NH(�8��r��Ҧ\�02������\��4Z��՟��G�0��[��L�ΪA���Ǹ��St��h�T�JDn ��a������-M�O��~�4ޓ���@l��l��n��=���#P�j2E�?΃xI��o�8��9�.�`L��k�5��ng��	T�J�1��씑�:��KY���sm- _Y���@�}%@�`�4��h�3��'c�,�[`�t�)
W�k��
�!���i��ċ�!-M�O��~Ӿ9�d�L�<��lԻ5�q�2��Kk:)���2�u]9�#�I�X��WG ���9�d�L�� *�P���Ga��T�rs�(�̴Y�{'%s�6F���y�q� ���+�6e���mn
V~$�zR���b��C����:�ɡ�3��-e�y��FlJ^d�d��l�v+�öJ|-���{1�����ը�k:)���2�%��짐b��, �k��9�d�L��s"�k
�5��)�rbJ6�~��J�����ը�k:)���2��N�g�c�` e8�~����h:h_Q\M� �]vAy*ط��wng��	T�w�&1�|���yG~F�Y��WwOkd��l�\a���5C�tTi���׏�����M�q�)]Q�x��r_��m�b�P�LƑϥ�g7U\a���5C�o<Z�L5q�j�r�(�EoO�؁o��L��j\%�	k�N�L�K�p��qԭ(K�l���`y��+a?��J�~�;��1��Z��M���5^sh�Qf�΃xI��o�n���� [��ѮT��~��׺���d�����G��Ð�gxM��R,ng��	T�rw�&�z<a��r�����?0K,��=���*� о��PW��B9�[�c��)�-9�4r��g2�~������\��4Z��՟��G�0��[�q�)]Q�x��r_��m�i��"u���Ȇb�L��B bb���H��efm�0z�cUL���ޤ�Y5x���:����S�>��a-6�Da�b�P�L��c�{rS�b�8Z���%\��o���h�Me!d��q杳/��-0��3t���=�4�04�jfw�&1�|���yG~F�Y��WwOkd��l�\a���5Cc�}���Fo|k�LbJ�1���K���L���4�04�jfx(�i��/R�*�W�Ǹ!2�͞nOY�c����gp��T=7�����bw��2V��K粞ƿ�Ս���:��֭�Q�>^��(�S�����O��KJDn ��a��[�~ē�J$s��(ko���Z��'��s�"J�CJ+T �o��_�R�wَVݳA*{�;h/�0h�5eש�y�k�A�$����@/��r ��9[��meF<i�LE� R8�k��z-�%��u�N�^X�!ހ�����|E�g�������(ӈ��Z��&61�~���i�x�0mo��[0�ʂ�j�Ï��	�Li4"�	��z��R��Y"�g�YZ6��HHD�u"�T�B�Z�R*E���&�Ut�\�@�\����@���kJ���af�iβ�=&��]
���b���M��#l/����1��X��WG ��<a�`�&� �EoO�؁o��L��jDY޶8�1�Z3�z:�������n2\�,h������v�}�@(H�o��΄x�g��	��S8�>���r8j�g����PTse��ͳ[�%�z�J���h:h_Q\o�HT蔊�cٰ�Ž��v�}����6S ��x���'RFtx�W��L�rw�&�z<a��r����5ߧE4��p�-a�D͢fU�9�׏�����MFi��|ր���5V��	��yx�_uE���З�Df�H��3�L�N ��HE����P�M��J{�����qθ�)�A�������>�X���D�gZ�w&�d�I�_Lm����1Eu��P�6y�J����+���C��엫��RH[�3�s1����*�|v�|-J�g]���V�|�^���X���鰄;Sn;�i� �uC��1Vhs�`�1�O�u���(%�9QD�Pj�?n�3��ϓ�g�I�*MT�*��\���?��9)�F��Q�������D{+�>���3�G��( ,n/XE�{+;3&wӱ-���R�t����ʵ���$�Ƣ�/�J�w��|��1�29tX���ʵ���q���� $���{?tQ#���<0�U\�BJY��~���0����؈<�Ҧ+��U���J����+���C���ϝ�HX&ci�=hkrHo�??v�x�[a�в����n�q�^ƩW?�d���&���m!q��]�г9�=Q�|?�T�U)��4Ps_*�GqW�w��fD4^y@�c;T=0��:ƥ0����%���N�s��T��[C��ԭ��20`��WV�#aطR
�^0oߙ�(ml���d����=z��k�8]o/�� �T^��a�@�nx���:�owђN�~u*w�A�c����sL]~ц	U#�&|R�� r�l6��_.����q�is���IX0F�M��LV�!��o�½X5�g�0�u�R'cf����(-ЀU�D�� �����A�{2pn��gn|�P� &G�N�g�c�`l����d���=|%��v����a�z6�F�KD�Vr[?z%CS2b-M�O��~�Ѩ�f?�R�:��er?G��g��ǻ�J���G�&&�����@/��r ����z�/���:����嫋�T�@�.��KT��Ҕ�5Ɇܾ�]��	He$(�2�ft+�f�;�>)�;��e~]1bt�Z��P��3�Q#� :a�	�+4D@&����1�qSm�G۞h�G�e�ԑ\�#l/����1��X��WG ��Ѩ�f?�R�Ԍ��Ǐ�c���w�I�7['D�C�k�a�	�+4D@i�a�sir
>Rf�����v�}������Ja�vݝh�c�A�L'B��o彍/Üy�a
��ү�+ҋvE7�MW�+�Dd�,�alֶ5mL�#���+�9-�i"'���Xw�j�7����	=��h��h���LX��WG ���]�UQ��D�gZ�w{�R�$�V��o{��:���m4��0�g�F}kQ1��xȀ��D�[b%Ɨ�tl��(Ur,J��`�om�c�Z�~c�}���Fo|k�LbJ�1��슀.�[ ٓ��so�-c�,�[`����_�=7�}|��	��a-6�Dak��"�՗�Cߋp{T���[�2�S�o��VH� p�;H2��I�
�2�j�ڴ���a�	�+4D@vE7�MW]��9��6���ʵ������v�Z鎬�������(�����?�cc��L=X�� �-M�O��~�r�^�#v��.ȅ��J���B�:����}7�������\�2���.Z��'#P�j2E�?��˓#���l����d���=|%��v��3t���=�4�04�jfrw�&�z<a�4�ڈt׏�����MJ�1���۪	�}a��[�.K3�$�)�vxg?�1xlC;W��A�eg�P�z��뜴����_6��&f<]jV��WD���Z@�����JYNd�l��?^�/k�i	��O[H5�Nw�$�^�Q�o�>�������7�D�;E��{oʃhh��;�H���oU�4{��F	�L�C���e����-���S�w҄ھɲo�I�xg�~p!ۓE�����y_�'�&r�Å��9�1|�Ҡ�ƆMk�	�X��ȅ�f5�5��x�,����L`z��KK0�RS�]
���b0�9y�+ð��T[�^�2�f'�^����t���3�l�K*�!b7�)���HŹn�軑��r���/�ciJ�0�I���!2t�ch������N��۞h�G��6�mp�#��1��X��WG ��Ѩ�f?�R�Ԍ��Ǐ�c���w�I�7['D�C�k�a�	�+4D@h�Qf��lW��ڻwR\�"mWx�W��L��w�򪥃WT
Y��%r_�1�J��]LB������([��}qn
V~$B�R���>_�zR���b�I�Q!9�{�����[�{7�G�7%u֛��B���EN��C�����w:qPL�
�*��_?�v�vE7�MW]��9��6���ʵ������v�Z鎬�������(����ЊҼ�<��L=X�� �-M�O��~���L�ΪA�%�C�5�ɇ����>�b��O������1�N�g�c�` e8�~���lW��ڻw�;����<W�1�.���h�Qf��&�(5�;2x���'RFt�T��,���}��֏i�RmHX���Azl>X��WG ��J��}0�^��3-����m]jx]�6k���cz�X
3kZ��\�G����s"�k
�5��)�rbJ6�~��J�{u(#��1	-Pvi b��a-6�Da�4�!���H�N��y�1�R�k�y��m�0>je`��@d:�����{~�;�z�G_����\�f�MX�xIh�Qf��5ߧE4������m����k���# m>���^!� wٻKm�Xn�
c����^eJ7�q���gҽd6U���b�%�C�5��#���H�Nb�*Z鎬�������(���4p���eqq� ���+�6e���mn
V~$�"L?��ٗ���#XNuK[~�H��1�>��mT~1�����(��(����ʵ���ه� �4�<J�1��씑�:��KY׏�����Mrw�&�z<aSm�6��`4�04�jf��ܐ�}�S��/:+�e6j�"Hs-�~A#ն�C;W��A�e��q�O�:<�..�4���Jk�����T��.���� s��?-+��퍜=jI�q|	����hV)_��s�֙Bb���dMA
��?�q�is��g?	��o�G���k۞h�G�q���01`��������ɐ�>8�co�v[�(!쥭*����	�������`|"l L�BV�����v�ـщ�l/g������g��Iw8�}�����>�EWz��ٴ���ad_t�5����3�����Qbݙ�-M�O��~Ӕ4�!���=�<�^�\�G���f^�V��?z%CS2b-M�O��~�Ѩ�f?�R�:��er?G�Wq�`ASβ�=&��]
���bιtQ�#��R*E���&�Ut�\�ً���N��A��J�E���V'/��������r"�F�*oX��WG ��)��]ӈ[x|h��8�iE�ı���Hҟ��\�G�����z 7	B���Si��i�
W� ���Pp��2�nw�q�u������q�k(��WV������'>D���E{��Ut�\�����F��Cߋp{T���[�2�|�P� &G�N�g�c�` e8�~���lW��ڻwR\�"mWx�W��L�7���n�f�hj�"��4^��)�d+������1��X��WG �����pP�h�Qf��n��K����P��+7��]�����V磆�._�g��%X=����X�3���L=l���[��Z�qѨ�f?�R���%\��o.��p*����H��efm�0z�cUL���ޤ�Y5x���:����S�>��a-6�DaѨ�f?�R�x���'RFt�T��,���}��֏i�J'l�z���n
V~$J��}0�^�s��R������f��go�4vu�݀�tTi����2Y��+rB�0j�䴑f��6�k�*x$6����BC?T��1摕\n
V~$J��}0�^��3-����m]jx]�6k���cz�X
3kZ���a�z6�%�C�5�ɇ����>�b��O����U6P�H�rv��qUt�\���	�Zo��F��hd���x4�#��p�ɟ�V e8�~����˓#���J��}0�^�s��R�����jv�'x�W��L�c�}���Fo|k�Lb���Sb�?�.oȈt�{�����[�{7�G�7^4�d'��{�}��ɣ@�[,E`th�Qf��Kf
�f� *�P����j�1>�+�9-�i"'���Xw�j�7��#�@(14~�����-/J�����Ut�\��"L?��� e8�~���o�z��T�t�x6�� [��ѮT��~��׺���d���ġ�j� |�p�-a�D͢q��`�LJ�1��씑�:��KY�[b%Ɨ��;�z�G_����\�f�MX�xI�P�HS|�4�04�jf�\�G���:��er?G����Oam�i��ċ�!-M�O��~�)��]ӈ캧xӍ.�-�f9@�~��O���f��J�1����ݾ-/�uu��ڿ$�)�vxe�zA��;��|B"�޾8�����q�]��ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0- ��Ckӏ�^!�:�_c�~:i��p�7��Z鎬������~/[�dw.2�҇�L�Xڈ*-È���*+��r�1��'p�@�̎�)6Opώ�,*y�#��_8\/Hi����s��.,����|#^�Vnl0��F��j �i7�sp>����S �=�[T�)��U�{'�$��'n�^0o����y�]@���U@���:��F�j{n�}�R �i7�sp>k�$����v7�'b����������5	��]�!���/H�5$�΁�a�n���o��C!T*�q���U�4_�;��	�'v�]��7G#+�Ǘ0z�cULOE��
����O�q�V���p��Nu�5=�����e�K)b��X �<z�q�,+	�q�P ڨ��S���Q�V�ɶ�w�H&���'ʢi�g�tpzl��a�|� ����7s�9���o��S8�����D�J��5j��i͠Z��)2��H�R�?�ˇ�h��<�W�.�P��:��Fy���H^5ʱle�~\3��Y�{'%sgeߪ�{(�%�8���0�W:h�o	�%�[�"ٌ�{m��ߏ�˯�h"E&��� ������`F�x >UZ�I�����w)КI���᮫J5�Hq�o�d@-[�v:v�o���+���5���L����;j�Mbѽg\��+"�9���B�I:׷�F�20)�_¿Y5��mn������Y�
�@���.*;È:�-1���{0Yaf�fL�!�]�BƠ���W,x��k8�5�>�yKYQs��[�|�F��˱4���[�jDG|��o"� ���I��Q�yt�G�^����]S�WI�;�_�	�t쩖NUD60L����L�Y&#t����n�~����p��l�n�Zlmך҉ݨ&@)�F� ��FZ���;D8���:��M�S�ᳰ��X�z���t���Xo޲G�����$7x�c >��}f]���]�w9"x�g�Hz���MN����!I/�������A��1��+�W�Ń�I��-Nd~�����)��ݱ�Ʀ�4������6�o8:4���8����t(&�L�\���F�`y6\�4�@���(�?<n
V~$�
�p\,%�M�_0-'h���>�,�V��j�3���!�`�(i3!�`�(i3!�`�(i3�it� B�a�a���v0�����c��.�a�9%>$I��h\9�G�2�d|�
�p\,%�i�X'H!�`�(i3rz��G�{0_�EA�������&���ΩL�*�1�L�:J��(�e,thS�c��}ZG{��7UZ$I��h\�oC��1_���l/ǋH��L�}t��T�s�)];I���8��/��o--ub �'�3�������r��)�=&�J�e�!�`�(i3!�`�(i3�����L�	�U��x]�i���E�< A^�XI�0�����&z��� ��=��Ɣ�S�h��ʺe��lf)��G`HE��R�km��K�Iɘǽ�������[�Iɘǽ�z� �����U�|/r��ऑ�y����Y�H~ XL@3~��k�f�U�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���aR���20�OU�	�|��><������p8�V�'�����v��K�7�wtMMC�)��3���]�я=�i���!�`�(i3!�`�(i3�g/t��5�Y�n!�ƪU�\HU��O�'d=�nϵu��3�5�����g��ǻ�J(��۝} !�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�it� B��~��ɳ�GV��)�m�g��ǻ�JƔ�S�h��ʺe��lf$���7O�R�km��K�jZ`��,������[ɨ�J���m
ɺ���!�`�(i3!�`�(i3��Y�H~ XL@3~�����Q_K�WL��<z2���؛y+��:�"��v}�\�����c�'��D��g��ǻ�JE��u1 )u!�`�(i3!�`�(i3!�`�(i3RN�]�5'�b1]�Q:~n�s~��20�OU���e�'�����p]��ܺN�K4,��Q7�wtMML��<z2��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g/t��5�e���!
�����_�X��D�VV}>iuLUX�Ϊ5����f��x�9�E��u1 )u!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�it� B��@֗�0
�16�l \�o��Ow;t4Ɣ�S�h��ʺe��lfL��<z2���R�km��Kɨ�J���m
ɺ���!�`�(i3!�`�(i3!�`�(i3!�`�(i3nTxꅗ�~�K^M ��k�f�U�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���aR���20�OU�y!���5�����p�~����cж #���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g/t��5�Y�n!�ƪU�\HU��O�'d=��K�G�5�������Oam�(��۝} !�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�it� B��~��ɳ�GV��)�m���Oam�Ɣ�S�h��ʺe��lf5�*G*B��R�km��K�jZ`��,�^$�cJɨ�J���շ��6yv!�`�(i3!�`�(i3��Y�H~ XL@3~�����Q_K�W�A���n_��؛y+��:�"��0Y��h�-��c�'��D����Oam�E��u1 )u!�`�(i3!�`�(i3!�`�(i3RN�]�5'�b1]�Q:~n�s~��20�OU�P7�?�䰱�����p]��ܺz� ����7�wtMM�A���n_�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�g/t��5�e���!
�����_�X��D�VV}>��6��J�5����̖�K �E��u1 )u!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�it� B��@֗�0
�16�l \�#����z�Ɣ�S�h��ʺe��lf�A���n_��R�km��Kɨ�J���շ��6yv!�`�(i3!�`�(i3!�`�(i3!�`�(i3nTxꅗ�~�K^M ��۪	�}a�]�w%�oφ��<�6���"�$�zf���&��7��������j4̗��W;��"r뾃	��s�G���[��N�+~*!�����]dKH��]�w9"x�g�Hz�k�>ur<&�+K���nC x�7*t�ͦ�J {s/� ���f�;�>)���K��<�Iz#1�<Td��"X��[硙�t�\�:��F�ā��O�q�V���p�x�*aE��w�����?OI�