��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-@���rahZ����*����Aڄ��[�k�|��ў��q����_�F��LF ��F9�>�^��M��7�m���<f#�}N9�h��/���b�%`F���\Zx�8��E��v�w��)?�� ! ,��e��~(l꼁��z��I._�O�
.�Zk�g�[��j�]�����8ɳ������F�A�xs̻��N��H^!�Kl�m�+�6��*��1�v����o�T
u�/%�O�"�F��� ��`p\x[���!�`�(i3W0�`��Ѣ�'t���/�!���c���"��z��"�����P��G�-�M��k�R��?xA4��^�y������9J�4Dvor0����.�q/�{<�x�fr��c�ZKY���#Ь�����Њ<s 2���ڠns6��������-VL�ސ���ƣ�L�/�\��9��IY���MTF�O;.��{C��|^����Yt��Z�M*q�M�/�-dOrS��E�����������I �x�r:�㜦��F?��߫�-H�/��� a�ik��Wʔ-�Y=.�"�K����X��֑xGV�M��T�t���(�zK�X饿��!��v����oX�$Z-�*��E��@��+'}���5M�YYroEێJR�VÀC�A��o��xȋ�l#ž��h�/,��ۿ����r�m�mIH3:Zt%��m&<�����9G�Ds|r�2?�����҃�F�� c��(�U�=��TA���#mԃw��+M}����j�����������d ���ѡ=�����Y �\Yy��V)�.�6C���Fz�k�좏1Y�_�R�|t�_=���$ۓ�����|Ǐ:�ues���$q��mKx"E&��� ��l$���D��Lh�Ԫ�u#7zǾIZ�Wl��>�;6W����F-P�u��.tƹy<c![���=$$h�8C& a�bD�G���O%���a\Y�����ḓ���X�,4�?n�[$��Q��3�O�2���Ė�� �Ueۡ萓'�al��p9�W�H{�G����g.Q�Q�?uG�)K|e�P4��&`��z��`5|⡰����r!�~WiZ��@Ő��thw��2r��h���\h��*�����g]��u�H1և���Bw��*`�|��K�z��}	�ʥ���S~:�:��3���C�P������eZ���(�Ow��/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'���?���ʢS����E@�ޗ9(����	�^��i���Ӿ���2���عf#�}N9�h�C����Y�q/L"t|Y�f�sJ�F���s�V�����<o�nïi�q{�f��a�:&�>��s���� T�8m��U}�	=�C��a���\�vūx`��:�r�^K������О.<�Ȭzn�w�'n�^0o����y�]��ӳ�Y�
Z�J
_�ʆ�In��tCF���y7�j�2\�{U�x���hA�4I^J<��H��&�ګvA���P`�|��K�zփZ���0�jݭ�F���h����tL���+��g�ڧZ��7�U�q��&�'n�^0of�`�(x���.j�,�3*������|���kJ_3#ڸZ鎬������rٮ�vF~�IK���Ig`i�ҋX����@�ڗe'���C1zh/�s��^a�T�~P�]k�!n}y���q���U�W����c�ZM�����{l�f|��rs�i�������k1T��v�܈�BT�^��a(􆿳�z��0������*�E��M@3%�w����$ĄҋX����`H���������h=-��;��lz������6�vg;Je'���Xw�j�7���|��{�r�\	��rR�^�V]��}R�wX�շ�R�������X��֑xGV�>�,2���7G#+�Ǘ0z�cUL�JJ�4(o�a\Y�����BT�^��a(􆿳��[ihC���%�ɏ�X,���֑xGV֚�X��M�TD���rs�i�>�Ca��?�o>�E]�٩��7�v�ԯ�`�L�i�C6�=�����!���;����J��6�vg;Je'���Xwb��Hg���'�r��'q�r.��c9�6�vg;Je'���Xw���e�KL[�#����KW�*�	S۱��J��q�P ڨ��S���Q�V�ɶ�w��V�k�j��ugM$BX���[��e��I�p\�WB�*�d��[� J���k�?�z7���%]��g���nU��X|Qeu��<�q{�f��a��\/�V����7�i���K�f�
�`�*%0�U�L�#_��^�+�J��;ۂ��IÙ=�HL'�kXyig@�����t��y�|�qx�]�V��v��K.Ū�C���D��j�69�$7��I[�x�]�V��v��K.Ū�C���D��^W�3B7��I[�x�]�V��v��K.Ū�C���DvW� �H`T7��I[�x�]�V��v��K.Ū�C���D�ӗ>���	7*6i��l!1�9���9M��I�� '����1��L��TZ����3;֍��@=;U�5V�˅|��k����z�KdL��[B�����؅��FJ��o�C���j��Ǌ�C��q�����/�~u+hBn�Y?v�<�!n}y��Y�{'%s�rOw������y$[|���"X��[z���6��+�x���+�qbp@���=ީa)��Ig`i�ҋX����f̲Az��%f�rE�X�e��Ig`i�ҋX����L$�����/���Ŋ�Ӑp�Dtq��Ig`i�ҋX����L$�����/���Ŋ��t��͝�u���Ig`i�ҋX����L$�����/���Ŋ����]D��;�č�Y���S�)37J*u�,�JL��ޅǐL�T�z�d6���|�_3#ڸZ鎬����Ĺ#{��	_1:Є8�Q;�m���!n}y��p�VU��Jm�QA�Q* �2��5���3(~s)tK��{l�f|��:2QYeƈ|���
p��v��֭��Ig`i�ҋX����L$�����/�Mv!���xl`�݃�|��].��'���Xw�����C�B�n}x��&�������{l�f|��:2QYeƈ�=�<�^\�c*�=|�WT�j
�I��w��,�,�JL���o:ϓ�gM��7P��T��TD���rs�i��ZIp����M�O��6a(􆿳� w�6p�d�H9M\��e���S��L�|[8�6�%ˮ�m�x���� ���S��S��6��o���+�@{fT�U�L�#_���29a���Q;5B5Y+�Y��d庒�D83��|��Yr���˩���.|�A6�E���?�.aݑMf���9���U� ���_j0��.@.�.H9���e#�|r�Mf���9���U� ���_j0��.@.�.H9���j��
�Mf���9���U� ���_j0��.@.�.H9��("�4��i�=�@��[�^������̇ki�D����m޴��eh�T�� �����r��T�,�'+���c[�u���褻��_j���=���a���Ѐ�uw�@.G5O7� ���Jg�C>��č�Y���S�)37J*uc�A�L'��-�S(�_Ma�~�Ǔ8���/�zeU�D�W�MԲ�����{l�f|�ό���.�܉��n* �w�-}�<��z��}�<ͧ�:|K5�w�x��?�����Ig`i�ҋX����L$�����/l◈�,��K.,�v�~������]�!���\B��V���)�xm���NX�c�|��].��'���Xw�����C����q
�o-x��az�d*�!n}y��p�VU��Jm�QA�Q* ���$þ�č�Y���S�)37J*u�,�JL��ޅǐL�T�z�_Flzk��_3#ڸZ鎬����Ĺ#{���0Q���ќבa��@IE�U����S8�	�Ms��3�˷���T�\ �������>�F����U���>$o?~�8r�k�K%*$�N�,�вԺL�9�d�e?��>ڃ(1����L�Y&
��L�>��ϣ'm�e��N(I:\����N��y]�u|�1��?��9O�������H��Y�{'%s�O��W��[�$��X�l�Lɼ�,0=]^	�&������%*$�N�,� :�:���H��߬���_;@�M�~��"����Y��ף��:����DZ���)i9%� MjC�9����T����X��֑xGV�}y���]D�]�!��	Ǹ�y85�}�-���O��g���ޔ�h���o�8���/�Yum�IʝQ�`)��kѶ���� 7⸠z�V[���>(��+ �\Yy��x�@eӎ��'������;b&��E���L��v�я̛��q������ �4���q���U�pzl��a��Y&��Y����C1zhg�����g��=Y��_Q2�+�YɢX�B���y%�ɏ�X,���֑xGV�U�(f�Z��L�4?@�T�q���U��s��d�\Hq�o�d@-[�v:v�o���+���5���L����;j����>^���o���KEd��]^X0��
x-	���'�$HgL��)�J����f5i�A��I`��=J'����r
���I}}3M�C,����|#^�Vn����o[���=^��>D�c�lQ�����+�7끍J�[T�)��
�6���.�֌���<�a)�m�d�so�}a�C�ub;�;��V�k�j��ugM$BX;Ά\C��ɧ���7�)a���%}D������h�br���lpda���\��6m��B��${��?�J�Z��]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gV��Vv;�Oe�d�#���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂f#�}N9�h�C���ߠ���Y��EMܓ���;�e >���l�n�Zlmך҉ݨ&@)�F� �@� ��LIM���zɦ�3y
�*����zEK#�E��Ǵk�?H�$�IX[��O2<������ #M�)��u��`�|�&�#�E�d��������y��Ld_���1[���K��&�|�G�2I�wp(��C�712��}ǞK=<^��`Y�F�����I��#��
Mcu�T�M�ڤ [�f!�)�X�j(�� ����n�
_��q���<�{�!���"�ֱ��R8v��j.Z��$�sӢ�]3�����c��(r$����GQ�A�����v1a{J���p���T�O
v���=�Ģ�U-��qs�VY��#M���N_��s�֙C�T&L�P ˃������H��߬������g�5���`JX׽oZ�j}�ܓ�s�8v��:M�'����f�����X�G[ᱽәBe!^p��X��ئ,\ަ�It�_���U�L�#_���29a���QB�P�[1�a\Y�����y�j\�c�V%q�9"�L�S��y^'R/	��x�◊n����E��̊�R�@Q��oL젡Iw�	::W��;1?�[F�9��G:([�(�����p߷T~ж� ��%lsσw�kzl`�݃�Tb\���~�IK�v���YI�L9@Ա���B������J�����P�'5%MY(璪��迿��!�6~[��M̤�1�G�Qc�Q�ޚ�e���62����^�i��e�`(\�ЕB;������E��@����U�p�6j�"Hsw��	Cʔ@� V�I`[���T�Յ��E���E9�Pt:> :�:������r�{"��1B�:ͫ��PK7'�r��'qm�±��m|� h�H�-�'�r��'qm�±��m|yʥb�9ɮ�c��W�Ч��7
T�%/���U� D,2(�a���g�|R��qH_��eE�(�������D'ڂ�+t�T�/7H~6a���u���i��g�7X�x�C��Jz*֢����X�M5���ʋ�1�?Ԅa�������:��}s��3�!�R�l����/����3��gL���'���[ЉiF0:��X���������̃��Y�����S�.�a����h�g���ޔ�Ѐ�ʲD;��|B� N,�N�'�r��'q#�� �[N0U�j!
�&kAע����X>j�V�����=�<�^����,�ǰ	M,��rER,-ڥ��-St��I=����)ڑ갚W�7E��,@�,-ڥ��-St��I=����)ڑ�$�ߪ;��hy&��-`�|��K�zµ��da��WV�#a��mJd��փ�G�#�j�!?!@e�کUCҔ[;H��B�O>q�j�s�t$�:�r�@Qw�c4~Nrg�d�/Ώ���я̛��q����#���/�g�f;[���e��@�Q6vmI/5(Q�g�+%f���at�)��d��X��WG �����9����я̛��q�����< ��x�-M�O��~�wq��Ǳ��<�?����k]m���ͮ;H��x�ԉ�>�5ߧE4��rw�&�z<a��N� φ��<�6�I���ftr���XQ �Kk�2��Z��%v�Ӫ(���/��m�±��m|4??-���/�q�Vٓ��(��������B}�%&^�nƒg�|R��q�B��S�,s�я̛��q����$x��7Lbq}��<�(���/��m�±��m|�c�ի�(_c�&��ʞ�sB�_̄�ѭ���m�Z9a\��8@0]�¯ץᝇ6H�����^�!Όg&W�w��fD���l׳d4��q���U�h+����~��Hp�J�,���tD2�����Vc2�����Vc2�����Vc��Y7��hx��W̚��j�l�����y�8T��3�u�l2�����Vc2�����Vc2�����Vc�-�������~ʪ���ց��_�4�'�al��p��M�.�͖'�al��/刲�Z�H���2	A�����e���X��֑xGV�}�q]A��G�s�� Ť�42��V6��xQ��g�|R��q^�s��Edv]̡<���\x&AAJ<�.6RV�������Yw�ōN����)�+`hBʆ[�$��X����$�PR�@��WPi��49\~���Y��,��9���	��%]�@�}���!���L3-�m�gib�U4ծ8\fZ�0uy&�Zz�I����g�|R��q��.N;R���U0��U�N�mQ]��P�$�����K��G����
��0��pS�I<�Y�Ǖ%�[.L�D�-��V�RDFR7�t�B
�6o�8��A�H� E4��/X	�HѾ�Ě�Z�(Lw��2?�.�����u��k�`���D�탯;\߰��&�՚���A�,�^�^���ԉ@0ӸQ/��^����c?��FT��~��)]��E��5xM�����?��9)K�C��m���*|�Ղ�];9�O���o��S��l��e1ێ�N�JZ�.�\Om�Z9a\��;z;�rԤS�
7�5@���-����U|��|�Tņ�8}��v�F#�5�~����p)'��:�Jlto��h�TtS�j��8�ɬc��WNp�m~|�ֶ��*��8K�ڠez���L�	��Q�xa��@�`��o'�#��A�]��h���/r�|��X���B�ݔ�]<����c�@�*����R����68��O/��G��-^/8��	��(Ks��0M�Bs7z�� 6�:}#�����@�>C �@nk�d�N�mb�"�i>8#��o30�@C̑<l��A�?J�_��d��N3�.���
�N$��k�(��Zx(j���q���U�h+���U[�t'8mQ.ZVRѿUJ�b��nw;��q�^ƩW?�d���&����3'�L��1�G�Qc�k]m��`_���U�u�!�(q��૦�6j�"Hs���O�ЉiF0:��X������G�z8����?��0SߖP�s�a&�Ep���f� 2dF.F?�o>��&{�'Y£V�F�P�_����3,�0/zﴚ�:�L��!�~���O�XA��uJ�9�ӧK�N:?y�gc��}	Vӯ)Æ��0��T��9q�b��|j�(b+���<�F�ۏn������F0E����țV���>ߜ��mN�p�b��D�RaQe-C��ʼ\��M��ڇ�e��M��:�V[A:�^a��]��d7Ud��A?Љ'�-�)0;S���:=�Dl?7^7]fn�c՝_�\�Zr�D�c��Qԣ��3��pg,lY����,l���8��g���ޔ$��Չ��׭!7y�x�}�0�.�,B{9��]��|M���/s5K��������K�}i�e]y]�g��i
E�ₔY	��W�UCҔ[;H'�)��@�D4�ky�h���R��%�ɏ�X,���֑xGV�U�(f�Zȿ䡜:[��;��s\ڽS�����4�֧��Le\`�?g��X̖�!=�MgT�����������h4c�b�md��:�L����E��@]٣�2e�tV��	��y ��f"���p���T������A�]���;��9�GKP�2�����Vc2�����Vc2�����VcFX��Go(�]R��w���5�5�_�vԡ3ѻ(ZH4~��2�����Vc2�����Vc2�����VcSd�*-}Q�#g��{����!d݊ܔ��$�����:�JH_�v�s�t��EH�a��㴺J8�����F,Z)����D
_oR���7@��-؞��i4��TH�a3k��\�'\��C��F���d`y���[a�^���Z�M*	aF�o�UI �F����X��֑xGV�05 S�s�l���X��֑xGVֿ!M�1#�Rr������;�' �2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc$��+�{c"G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F~�?|�[_wȵ�e�kY��Y+]��=W�֯�^��N�&��)��m��[4�l��r����#�[�+��D1t&�B�j�O��(a�&�<��˰���,U��2�>D�c�lQKݗZ:���'n�^0o����y�]�'�3�$ �#^�Vn�^ֻ����XP��ȭ����m�cc�PƐt
׫�J��q{�f��a�:&�>��s��>��!���t~'�^ֻ����XP���a�=U���O�[�$��X�R>Gn�
�;5B5Y+�+�����E����z��2U\���\8�ǔ4�_a�CK�H��=�e\gn��_�G��G;5B5Y+�T�����N�a-�E�S��i=���[&��?��
q{�f��a��4�6�t� �R���({&3�-��_�s*)F����'n�^0of�`�(x���.j�,�3*	��<���u���d��CE�-�EU��P�:^�J�_-�_3#ڸZ鎬�����%�����~u<ѥ�"���$v�~������]�!�����#e;7mg�oc�.[K��m��/��*(�I�y.͸|��].��'���XwZ�֢t��FC5��v�c�.[K��m�u�M$S�{�,��TG���|���Aɘ%�ָkd�vu�Z��F����{l�f|�ό���.�2��T
�r��<Н?b���-(S�)37J*u���
6��!l$P�ĝ�����-�$�<��z��}�Q2�+�Y��0]���!Vf����aU�7L�<��z��}拋ġC��ױ����h=�R��a:߻�%�q��{l�f|��rs�i���ZS��0���@	Q��"X��[?�e`N�a�� л��{ET�\�%�OǱq�d�ֳ$7bOc� LҪ̆`K��"ݱDˀxRH�_Jz����I�����KW�*�	S��@Ő��t���N�kcI��S}H-��;��lz�������{l�f|��rs�i�>�Ca��?�o>�E]�٩��7�v�ԯ�`�L�i�!s"֛
.C���~���J�������L�'���Xw�j�7���|��{�r�\	��rR�^�V]��}R�wX��0���7�0>�Q�k^�ïw��O�$F�|��].��'���Xw�c��Ut�#mԃw���k]m��8k>6s����]�!��	Ǹ�y85�}�-���O��g���ޔ�h���o�8���/�4��ľ)T7�9���������D�7��S�:I��w��,2�r@ڸW��, #3���t���(�xIȀp/x���̝Ʃ��&���#�{�0;�}��Ls�����D1t&�B�j�O��G�Z�4{�%a�E�IO�#���O	f׿���'Y��6��X!�LHi�S�������GJHn��z���u\���e�^t���*��E�V��yd?s�Nmg%���ϯ�ad"��g��|���@!~�X����Ѵ���/z[f��ϯ�ad"��g��|���@!~�X����Ѵ����&����"dϯ�ad"��g��|���@!~�X����Ѵ����F.BT���Q�����aw���Ir^u%��ӻ�VH9��h�c�!�洵�q~Y�a4HSwk��m��\U�L�#_����Y7�Z�1�9���9M��C�0� 9��@f i#@���%&E����T�;��s\ڽ_3#ڸZ鎬�������(�����7$��t�Ȯ��ߊ�R�wX�ղ�=ީa)��Ig`i�ҋX����@�ڗe'slxSwP6�č�Y���S�)37J*u�,�JL��އ7m�~��5ч/��n�v�~������]�!���\B��V���)�xmB����B���|��].��'���Xw�����C�����d�W��!���{l�f|��:2QYeƈ|���
p��j�14b>���Ia�i<��z��}�<ͧ�:|f;[����[��B�_3#ڸZ鎬����Ĺ#{���g�.���/������!n}y��p�VU��Jm�QA�Q* 510*���8k>6s����]�!��	Ǹ�y85���Vԓ4��[Ø�;�x\�HP@�a����U�p��
���)��ZbMHmH�bȡ=s1'���S��L�|[8��<�yi�B}ْl��]�B�M:��2�n�ڤ����]���uc�_�����.dp������'|�?�<�d�:O��?+��9d?�3�7E�7�<��q{�f��a�:&�>��sU�L�#_��,Vit�-k�T[���e��؅��FJ��o�C���j0e>r��;�[qo��Oe[B�����؅��FJ��o�C���j0e>r��;����;-��[B�����؅��FJ��o�C���j0e>r��;�}������[B�����؅��FJ��o�C���j9Xi'�μ	����t�\x�]�V���\���Z�-ªQ�C�ӭ��n)�T�ژ�k��Mf���9���U� ���_j0��.@.���=��s��{`����!v" D��ﺣ��{l�f|��rs�i��ZIp����M�O��6a(􆿳�����?<��"��Uە��>����V;5�č�Y���S�)37J*u)T{6T'r_���#��v�~������]�!��5��E0����)�xm�v��C�xv�~������]�!��5��E0����)�xm�}�Z�t�v�~������]�!��5��E0����)�xm%��eG_3#ڸZ鎬����Ĺ#{��	_1:Є8�/������!n}y��p�VU��Jm�QA�Q* PㅇO݉Mn�(�At]�<��z��}�<ͧ�:|��u�읛#��Q5����Ig`i�ҋX����L$�����/l◈�,�!�1(n_v�~������]�!���\B��V��a���	�YI܁�條{l�f|��:2QYeƈ|���
p��"h�u)(��Ig`i�ҋX����L$�����/���Ŋ��\�c*�=|�WT�j
�I��w��,�,�JL���o:ϓ�gM��7P��T��TD���rs�i��ZIp����M�O��6a(􆿳� w�6p�d�H9M\��e���S��L�|[8�6�%ˮ�m�x���� �K̡g��b��M894��f׿���'Y��6��X!�LHi�S�������GJHn��z���u\���e�^t���*��E�V��yd?s�Nmg%���ϯ�ad"��g��|���@!~�X����Ѵ���/z[f��ϯ�ad"��g��|���@!~�X����Ѵ����&����"dϯ�ad"��g��|���@!~�X����Ѵ���/U���!-�iP��G��x�]�V���\���Z�o�C���j9Xi'�μ	����t�\x�]�V���\���Z�'F���t���s�ۦ�*��z�KdL��[B�����؅��FJ��o�C���j��Ǌ�C��q�����]����+g���wƱL<��z��}�0z�cULm�%������:F�X?�g��U-�ey) ��(��?<��"��Uە��>����V;5�č�Y���S�)37J*u)T{6T'�D4�ky�v�~������]�!��5��E0�u�K�]���=�7�V�_3#ڸZ鎬����=���ޒC>:G�b� ���Ia�i��-��%M�:2QYeƈ|���
p�c�+�%I���Ig`i�ҋX����L$�����/l◈�,� Q���/v�~������]�!���\B��V��a���	�YI܁�條{l�f|��:2QYeƈ|���
p��v��֭��Ig`i�ҋX����L$�����/l◈�,���ؽf�����9�dMbZ鎬�������(�����7$��t�Ȯ��ߊ�R�wX���"h#�)��*N/�p���(�
t�������2����U�p��
���)��ZbMHmH��R�Q��=O��'�>�*eg��:����H�6�
�Ф�kg��')Ri��뗬'��x��H/�/UMê�[��M��LG�IÙ=�H.ZVRѿUJ�b��nw;�J�l�u�Ã��*=M�cu�*�.u%������Z�M*�Fv?�S����0��7���Y��Kd��TGcL2���o�7P��T��]�!���o��w���Z7N�ש��*�U�t����wi��(S�qfm���u��Y'Gklʟ�����Z����d�٣�����6>���T~}���T>\��&��\�4����ﻋ-��Ȇ)��e\h��K�Q���lp��z��a7��ﻋ-���C�M��N�۔�Zr�lR�����i�㱩� ���d�٣��5*���ӡ��t������lSԃ���~�:\�h�]�!��	Ǹ�y85�������IeuѴ�8��ӳ�Y�
��m_�\���8���/�a'�<� \:h�������j�)䔫Sx�lޞ�ό���.���K�Q��L�
�T��i�Mf���9���q���U�KX�U~�?)tI3�;f�ӊ[�k��d�٣�����6>�����U�M���sp�	O����ެ@�o	�ﻋ-�����S8�6��s*3�$�Y
 ����6?L����[�Fc�k��`y���pzl��a��ʳ87��Q�
#>:����0^��V)�L:�焘q���U�pzl��a�K;���DG(K�Tl�;���f������=Y��_Q2�+�Y�����n9�{�]���q�GR�Sx�lޞ�ό���.���K�Qmd��gޗ� �4A( 6��D���Z'���Xwa'�<� \����9%=��M]l]�Qbi'D�ﻋ-���C�M��N���N��+�|�1��?�WdM4@Ȍ[PP�\��]�!��	Ǹ�y85�}�-���O��g���ޔ�h���o�8���/��6%j_�zHq�o�d@-[�v:v�o���+���5���L����;j����>^���o���KEd��]^X0��
x-	���'�$HgL��)�J����f5i�A��I`��=J'����r
���I}}3M�C,����|#^�Vn����o[���=^��>D�c�lQ�����+�7끍J�[T�)��
�6���.�֌���<�a)�m�d�so�}a�C�ub;�;��V�k�j��ugM$BX;Ά\C��ɧ���7�)a���%}D������h�br���lpda���\��6m��B��${��?�J�Z��]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gV��Vv;�Oe�d�#���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂f#�}N9�h�C���ߠ���Y��EMܓ���;�e >���l�n�Zlmך҉ݨ&@)�F� �@� ��LIM���zɦ�3y
�*����zEK#�E��Ǵk�?H�$�IX[��O2<������ #M�)��u��`�|�&�#�E�d��������y��Ld_���1[���K��&�|�G�2I�wp(��C�712��}ǞK=<^��`Y�F�����I��#��
Mcu�T�M�ڤ [�f!�)�X�j(�� ����n�
_��q���<�{�!���"�ֱ��R8v��j.Z��$�sӢ�]3�����c��(r"�o�Q�EZ{�^�#�ZeT����7�@�0�r���a�)Z,�9�GKP�2�����Vc2�����Vc2�����Vcj+�;H,�^��Q��+I�[���ca��&�&-�(ZH4~��2�����Vc2�����Vc2�����VcSd�*-}Q��kL=�F>��o����o�fon�_�(�8�"�~;ѥ�RKW�*�	S^�����&s��חo���^hY'm0���?*е�^���wƄ�{Ƨ\bT]��7ۺ�#�����~��l��1aΉ����ߚ�����}�A,�S|��4���dq�e$��ӳ�Y�
ۼ��	K���$�(�+�G(��Y�Vd�8��N��(��{̑6ԉCy�8j�Y����I�k�%E~���J��ҝ���O�B���\媠 �eqɟ�R��(Q�u�<�w�i���2XC$2/G1�ԠֱTU8-R�T���k����$�����K�ֽ*�e��J-�1�q��)��b�Q�G��-�siË�M{z�(�˷�p"�.����L1�%Ŗ��g��T�/���B^�!n����d_��s����I8ԗx f�g\��*���?��c��R�?��Xq_í�F�s-w�?��?h�F�UΘ���.\��g(4��4�S�.u
i*�TWT0z��~�(E�POlb��]q������WV�#a�}!Z<>��V��&|6�łZ��0yI�[	ϱϭ����y>��v����jht��g�����9�g�klʟ���Q��:'�TPs_*�Gq�p���xg����6�������C;����Es���F1xk�k���L݁#g�k��g?	��o^3�|J�܄��� M{��(:/�b�&�q��ث#*�	���vAb@/��r �>/�w-���V��&|6�łZ��0yI�[	ϱ�f;[���v����jht��g��倉r˲���[yfX��[b%Ɨ�^Zp����4��x:A4b��JB䶓�([��}qn
V~$��|�;�#klʟ������u�h1�@/��r ��%�z�J����C���Uȓ�z�������C��R*E���&�Ut�\�8�8��gv8(?i˸3�J�
�MɂMv!���xP�o��x*ȩ��>d���,f1P�y�B���2L��x�ԉ�>B�R���>_�{�Z՟|
[;T�!'ؔsy1�n��뾦�f ;h�Z�O�#��K��%r]�Bа���/��D��c�Z�~c�}���Fo|k�LbB�R���>_c�Zਧ�%z��"�����P��G�Q"���_ނMv!���x8�8��gv8(?i˸3�J�
�M�'٥��gV�J�1���K���L���4�04�jfx(�i��/R�*�W�Ǹ!2�͞nOY�c���1�ā�����-ĭ5�6_ �nޝ3���� ��ɔ������?���;�$Y$E�B٘�#g�k��5د�������f�����X�G[ᱽәBe!^p��X��ئ,\ަ�It�_���U�L�#_���29a���Q������<`�y�����Cn%�}AU�L�#_��^�+�J����������@	Qg�m>�`^���t��˳�M:��2�;�琾BT���h�}q���'U�	�YI܁��DCX�.C��1�gB�� o� c �d�N9N�510*���IxoҢbu�g��A�i�8�=w��ir肃r���4�磕shf(�`�X�G[��c�fm���3�%Uo�'�D��¹��g�0�u
��"�!�sp�	O�ƻ��W\D�F3���%Ff"�	-7���ү��d�<��7���n���&�Pݭ��%�x �ǤZb�`�y�������"�X���G�����:�5Ӡ�X���e��
Ut�\�5�UI1�gB�� ]�Q%�n��뾦��"L?���P�o��x*ȩ��>d���,f1P�y�B���2L��\n0�8�:䩒=]'���76S=f�?TY�ސ�����)G�J�cbp��'@
9��y��%��3��ןmnRYpW����@	Q�M��k\z�$Y�G_Q#j<��#���z4�����i=���[taT��bX��WG ��v����jht��g��倉r˲���[yfX��[b%Ɨ�m��"���@��b_їE����ݾ-/���b練5د������
#>:����0^�� ŷ�[�}Gz�F:�@"��]����ڙ�����r(H\�ܢ��,	սL��$����,�ǰ���[�F/$�J���3Dm��A���%'ף'������d�l�'�al��paf��pD��>tT��N-بS� �D���B]���L�����=4�&��Q(I��M@3%�	����,�czb^y0�, bާ�kU��sC���X�45إ��ZWuȅ��SZ�N����VM�d�ꂕ0.p/��sH�}ˮіs�����������,hg~W#_pCeu��|̙1ږ���[�$��X�aM0��x9@xi�n��\ؤ�z;��$v��g�>�;6W�e�9�s[�A���t��˳.D,����	�YI܁��X����{o��&��;��L�Bza��i�g����l�1�ԀU�k�L�Z9@�;{�����%����%9��T�ِmd���u�a��bZ1�C�O�hh���X ��Y�����Y'b�'=�(�Ō����,��5si|�1��?�WdM4@�Z���}h
�#mԃw���k]m��yʥb�9ɮ2�����Vc2�����Vc2�����Vcv�iL�D��u]%_�ل�����5IΫN}q�~#�\��V2�����Vc2�����Vc2�����Vc.�
͹U�M�C:4�ֈґ�y�x�Q��C�uS�4q�
t�DY��b8!�ì�	jM�C:4���"r�V����U����r��<Н<�Xo���$����?�܃^�Y1V�&�i�д �rH:F��
 {�L_k6�iUrx���p#�r6�x5�A,I�@�"|VD.�+���s�f�I�w�U��|���1?�g��VĚ�d�>I�~�щ�X~��`O�g�q	G�Q��q�ﲾ�Bە��'��e����9�����Q�b6��pB0�iY�<�C7F�=j������<Va����7.N�ӃHF��v_}M������}'�=�+!�"y�W��n�)��o'>���?����u;϶i6����R�KL���:� #F�E�Zgu�t�1g��X��ن�	�a�B�����3����L�Y&Kfȵ3�\=�r}�Wq�ꑉ�� �3��l��gS#�-�tS~1x0PAok��G��]_$A�õ�٭�����ґ�y�x�l<Gt���{�]���q�GR��'Sդ�!��_S1�����o�>�5�Ǜ��k����>�lIorǟD�uiM���	�fmt����]$�﹈�i�~�Ԣ��D{5���U�L�#_��,Vit�-kݔ�yN{-v\L��"��#nS#y����m�(�����p߷Td��#���~$�q����!��ZB����=�+K�������үf�D r�f��h�3(~s)tK�h�RZ9�Y`�ِ{o�7���B�=�7�V���үf�D=�
�a�� D��ﺣ�i��¹ ^��y}$�)`� ��qQ��R��-���fx�Z�0�ԋ�Ƭ�����D�� >r�Z	�Ia���F�笣�.Z;�������xa��rװ� t��]�qa]�݊3�m�E;���20ӠH��=w�A2ޮ}'�=��~6��_��jt0��Ƅ^�=�]�_Jz������D��ܒ0�=1E�Êp!!v*!��4�b�Eƃ��Q-s�b!��u���͂EC�y��Q28U�sQ��=d�Ɇ�X�$Z-�*�����-VL�z����9�j��f6&��?N����Sr� �A����ҹ��)U��XI��ׅy&�Zz�IÛ	���~��s��>�̔���c�(�3��[��\*n6�-�Ƙw���+t�a���`������w�=u�A��7X_��7��W`i�X�QK6�E����*��[�$��X�l�Lɼ���C�O�d�xǬa��u����9A���q�O�����¯�P��C	,��Ȃ�	�����'C`ø�X�t�G�����u�����&�܁�^����r
��Cݮ2�����sE���y1+�줥G��j�D�EH<J�B@��(�hS�}e�܍ˢO�bF_��a��Mz���O?�Sկw��[#M�4�!�["[:����!��lSԃ�0�!𨱹�I*�?��m�±��m|�Mpl�p�;�s�*�:�L�������-VL�++��Lm�>�Q�k^�ïw��O�$Fg�#辭aE߅'O�%�z2�^4�l���lp����0�Rݯz"��G���P�f���oH�pNM�M��K�t0�5�]ؗ���0�E>�z�>C��?\$��M��ݺ|��W�_�\�Zr�2��_:��y$[|�h���X �õ�Y���<�&4]��W�q}�w|�/U���!-�iP��G��\OL^��>%�Нo@���;1?�[F�sp֟kh�y��;��lMԲ���L��S-�����$þh���X �����R]Y�3�#�����T<�t�S�@�l��tt�G�d�d�+��b2������ȼ�4�!O7I�"h#�)���w%e�D�m	$�WI��)A�
��v����=�\[L�R�X��Uq2��Z^��:�C�7�]���GljJ���a�X�� ��v|�ˑ����p|3�f0{��
�� �:&��L&fL0