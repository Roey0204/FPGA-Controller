��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-Ǎ�x�"Ec6G̑�|̍Df�z�g�����#�=�[.>��$^���?�G�P�U��:����E;�i�:��ꄟ��;%�"&����XX�Q_f����N�=1��1��ʀd3��ş���L:�%����:}�8�(�2JF�E�bU��_#`k^D��ń�"&}*	T��(��gjq�=?ل�Q�g��6��ە�q�G@��LF�+,ߩ��A�^����*�^����A�F�7���3�GXS����E@��~���($�J.���
��'p�@��rB�6C�2��G�����#��%&�� ����q��>��yܛ�	��|��	(���zL͊�q����N�:�Pn���������W;5B5Y+� �i7�sp>7.~Ƨ����?2^�9<o�nïi�JHn��z��r9�3�X��-�`V-u9�`�jݭ�F�����K-psܧ6e���Vx�ӣ�3�9����Σ6��u�_����+����U��M��f	����[I����,Y[��FzBR)�5,F�ʦ!�_k�%w�_3#ڸZ鎬����Ǟ��݈�Z��l@+�v�~������]�!��	Ǹ�y85��r>?�W�p��HM�e��`y���9��
)���l�F~�h_3#ڸZ鎬�������(���}/A;T�c�owђN�~R�wX�աzZru.��'���'X��6�vg;Je'���Xw��%�r �&M��y��Iۊ��8���K(��z�j�;9�e����E�$��1v=��`x�~�I+�?T�]D�9�ϑ��[�֖�9x��i��&��TD�Y�J7��e<�1��bÌ�s��X�e���V!���IÙ=�H�^�p"ORmHX���׫�J��q{�f��a�:&�>��s����ӓ��^hq��:�}0�st&���\�v��Q���K�c���%��a�����*�����Ѣ�{l�f|�ό���.ӗ�!����jT%q�#�<��z��}�Q2�+�Y�slxSwP6��B5x�S<��z��}�Q2�+�Y�- 
�@
���C�����7G#+���[H��Q�$�k\_x���� ���J���_����A�2��G�
��吃1�ﻋ-���C�M��N��[XJ[]WQM-���G�yQ��Z鎬�������(���}/A;T�c�owђN�~R�wX�Շ��uj�*��MN����!I/�������A��X�@�5��6�l��s�����[� y�~��ż3���F����T�O�H'�J�����=<�HI����>�W�_=��0���̏�u�=Cm�v4��61��7a	�����Y�
ɸ�oƴd��t�'��9ܛ�	���V[�+
�l掝�K\m��U}�	|^�׽R�s�DH}�_z�9�E�\����8�i�`!31u��9x��i��&��TD��E-%Jn��ɧ���7�)a���%}D������h�br���lpda���\��6m��B��${��?�J�Z��]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gV��Vv;�Oe�d�#���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂��(%�9>��!E)ėתJ�#�P���(V�0r�����K�9y^6gV��Vv;�Oe�d�#�
�{�-�������@0k W�:��S��y9Ez��}��H֞��� �0\��.�g6���@�H	)pH!���5�Nn��XLVt����G��5�On"WW�p��G��8���Y�઩0g���>{@�w�|���*��>
�-�E��{���dʡ��'��gk=���G��yʼɊu�V&��F]�&��yJ�y'��BSz��w����s�%Ƥ�/���d}��[�ƭM��g������Hhqu!���5�Nn���4L"�+�va��2kYD����������~����MA�q�m�,&H�[&-nD�P�E6�k��q��־�h��z{�;r��E��Gή[*%��J{�+�M�( q�$dШQ;�im��|�L�݋rq�_���13�׍����V��ÑR HjlU5oܛ�	���G�˹Ď�֡�\�<7�X�e����]��m�n������"���P�3 Ei;r�.�/'�����WX�*�܁�c�PƐt
�G���خ�c@{���(f����zhc���>��3/������ї��*[UxG���0`K%Z�<�){:z��!��� �9�Q.��k�2��$cIn-Hznk��HDL|RIT��q�0 �_	2�;j�ٕP��P�*w.�S��rfz��	j����.�hXQ?D�BLM�s�mP6�Ee�&��c�����|�\;͖�"�Y�%u�8]-̧Z�hXQ?D�BF������l*O����v=��`x} �0�1�c�Z�~yq�Gw���Dq]\�����@	Q��[�Fc�k9���.:���B��U���-IH�"�k
d���I�z�$�!�a��o���!��(��M��|���!�6�0?�aV���p
v�ݾ-/�uu��ڿCt�w#��@�������a�U�ے
- 
�@
�_�-oH;�A�߹�+%C�@�׆p�9������ �ı�ZnZ�^6N���j/�(SB�� X*�R:||�T�w����]�*�1K,?�ƕ7�F~؅��'�u�u������k�Nfz�ǈ�,�Τ�D�w��[#M�E��Q�������'Y��a1�Z���t�K�"i��I�&Q�P�ۯ>�[��b!��u�,ҹ�$�d_����M��S�	RN&�����]qs�)�*6=�z��z���Tr�-:�����
���*,f$�7Q0- ��Ck�fÜ�2/�ri�y�!�3���1�/6���1@�,wLn������ْl��]�Bu�h�ɟ�B�I:׷�F׫�J��q{�f��a�:&�>��s���� T�8m��U}�	KݗZ:���'n�^0o����y�]@���U@���:��F���V!���IÙ=�H�swFy76�$t8[�*.%��W1�č�Y���S�)37J*u^�6:���heJ��Dv�~������]�!��j������9��v�~������]�!����^]����qZ�L�8k>6s����]�!����k>#%Q�q㧵�0�!7���kv Oag�qod�֓��Kl߯l�A�߹� ��F�I`>�YR��jG�D��:�3Ϛ�ҋ��Z鎬����Y�V��#q�G�����~�1*sukXԙvh�q���U�g����IX0F�M��ȳ�M�|���!�#�xd�< N��r*$7�门Q��Ȝx� uŤs��_ɇ� ڶN(���:�A+�\��N��-M�O��~��r�t�nI�w��[#M������Ut�\��V�.5�i�[+�bna%��w�G4�4��w��[#M�%��v���@u��B�|���!-3��MN�=�<�^���pP��G4�4��w��[#M�n��뾦��@u��B�|���!-3��MN�c�Z�~p�-a�D͢q��`�L��˓#�����V|>�b}A�<c2;�gWaU �I�%�z�J���'Mcö]�q9+t�}��"n�Κή[*%��JGjE���%��v��>je`��@d:�����{~�'Mcö]'�^������"n�Κή[*%��JGjE���n��뾦�c�}���Fo|k�Lbx(�i��/R2Z�<���tD|�u�@�A�߹v�;D�}�f;[���x(�i��/R$ty�h&������}-���ǯ3�4���4T_�wx��|�w��Q�U�k�
�^6N���	�<?��%y��Pw�54�����w�����?OI�