��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-~09h�i�Nq�{5�h��%��Xcbp��'����Q4KҲ��r�D� �m�'�t�חEʭ�3�Jld��q�G�~��Z2��˝1~OT������oPY̅���c�PƐt
׫�J��q{�f��a�:&�>��s�z+/�c�Z�J
_䆼�\�v�����{�{\J�yG����y��\�vť���ҧ`�S�*H������=t����w���@�|��].��'���Xwd�n]Nِ����_H;a(􆿳���A�b,�my$�N���Uە��GV��y�&_3#ڸZ鎬����D�OBp�b}��BB϶q��{l�f|�ό���.Ӳ�[O�"���Ig`i�ҋX����@�ڗe'��E4�Mʸ|��].��'���Xw�-X��-���Ig`i�ҋX����@�ڗe'�@.�>�ȼ�|��].��'���Xw����UA����Ig`i7G#+���[H�����2��~��o�b�x�'�6LE�EYZ/���)֨9 >�j��O0E>�������fHa��!A{�H]�%�Iߎn?�e"�2ao
r��FE���r#�9l$���޸�����C�O"I��MjX��k���`���F(ĕL2	X�vb�)�S�����]�c.��'1����1\���k�e1i��Q,�&d���ݚev3Y�IkT˱ ��O�������]�U�����8�o��@�<�qؚ��L�NG�>)�����7������7�� �����R=�;@R��Ω�dBj#/����@$˺/tw�ԝD=��٭@�FϟQ�-i�`�g``FD�e3>�ƙ�Ǘ���mC��XH�����wI�d��`���1�E��)֨9 E3����=E�EYZ/�@�L0�6#����"'W�9�p��y��9��L����Lo�I��'��恭�h�I��'�%�e���Ĕ^ֻ��X�x%}�����
D�5tm�c�oL�~j�F},M�5����`K�����svfY������;5B5Y+���o�(�)��;U��tm�c�oL�������FTVP��b�M:�8U(�d�٣��c�A�L'��y�!�;&����˚�T�\ �����j�|�z#:rQ��q�X�G[��;ۂ���cY�~�"���ʷ��1�(ʌ�N�M8�U����t��h~��J����^Mf���9���q���U�pzl��a��i��؂ۃ�y�wjאﻋ-�����S8�l��`�_gi�.�!����Wy����`y����s��d�\��MN����!I/�������A��X�@�5��6�l��sХ+�:R 8*!Ē\��c�PƐt
�20)�_�5�e��a)�m�d�so�}a�C�ub;�;���A���g?�뭨�fv8���p�lő�4�`�+��t�Y�Ij9���"]�ɋ|5���F��S���v�@�y�L*���8�^�.eO��q��S��;�(e)��v��=����'�$��u,��y�"���Չ-RW!�՗"<���^[ �1y�,	��"k@:G�	���=�ܾ�y�c��"x�O|?.����!��!����W�������9��~j5��Fo�P2}�).;��L�O#t����n��]ߺ�`@ZWH]�+�a�/��/J!�w:����v�=��Kܷ��=tʻT׼w�V��r�N���7B�Im���'��P��+BY��9���$�+���)q7p�5� %�����J_�xd��j��w�怖��CcO^Z}��"X��[�p C;8;�IX0F�M��2��h0�u< j0�l���zV����l�©T�rM�W˳͠m�xW��-#��k{-���#��H����E����d:Pe�KX��ik
>wS5�s�E^Q�-��<�zD���z-M�O��~Ӹ݊���K0�u< j0�9�դ��8-M�O��~���t�)�A�ސ���U4���Z�+�����Ur�7��霖�b�z'hۉ)��R��삠e��@���8ᶉ_x{^4��*m�D�$0䤥?��a�&qԲ���L�x{^4��*m�9�d�L�D��7��(���W\Dܕ�%�������&�����LS���W)��/807���>�V�^oa)5�(�� ���$�I��#�Z�����nc���m�vG���:�����"L?���BP{^�~m�(��k8�C+���Hm�(��k8;��_b(�c�}���Fo|k�LbS��_�ɤBtL+w�}��r��g},MM
��,={H�3)-.�qc��.�g3"F`}%Z/�Z���m(f�9���s���C����H��+��g&���Fm��Or%+�"ɽ�gW���"���甑�:��KYCt�w#��@&����1�R�S`��sK~���mv����͖n.�v�L#�?�-�Vb� �F�t0��0tm�c�oL�;U�Qb����ג��ryO#��!�Y��N��0��汣��~��#k�˟ܒ�o|k�Lb�5ߧE4��J�1���k_���b_!2�͞nOYA�	��7��i���]�tR���)֨9  ~�G�	9