��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-~09h�i�Nq�{5��]�0�lK'���Xw����Q4f����om2�YQ}�U�"g%�\�Ji��'��%�a�z�o���Ή�����f�p��G�42c�Ϡ\�)zL͊�q�� �^�ߏ'ER���c&;\e�L���'��-d�Ry��\�v���T�©ޒ�����s�VKOi�~�n�
���b����Y�{'%s4C>-��3v#��.X���*"v%)�����iR˳͠m�xW�g]����n(���˧[(X�#��§S6]Z���榡dB� L�s;X�a\�/���~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢS����E@�gh1���Yh�\��q,f$�7Q0- ��Ck�4���_z�k�۸�y�uZoO�=���t8� L�s;X�N�N���aC�h�>��!�̰���_8\/HiO���L�~h0%�������E3u�;5B5Y+��q	k���A�XWf^64W��^�o�A���,r�s��pK�����o���M��JVLM∓/^
wUgJ��Kʸϸ�N�
�o��djf[P�O�+`�W��� ѦV��7^�9 �;���b��iAj %�Ho�-[�v:v�o���+����7X��U�?	r���g�0�u�w��$C��׫�J�є^ֻ����XP���-O/ [р$	3�Ð�9�X�e�b��@�zL͊�q�����芶t���6��^hq��:�y���OJHn��z��r9�3ꓩ�l;��!I/�������A��1��+�W�Ń�I��-Nd���L��)�1��b���H;nvļ�\�v��	��2�Vz� �#'�a���z�&���O�ukQ����\{��x�gPo���}ђ{)8A��;ۂ��IÙ=�Hmn�}EGc���E1i���7��q�2$��\��@�n��3�op��м�\�v��&��DZ���� G��t1�.))b�#�\��@�n���c�SV�^ֻ����XP����j����@�w
��о��PW��4"ۓ�q���v�4FL7D�6�~z��KІ��������5�2`b+�\��^ֻ����XP���%���Nr�X�r���eC�!��6jV��������a�2�`��I��3+��96�ltN�C��NxU�^� d�Ew�S��u�naJ1��\�vŹ��7���J{+�ę�^�"�S��_:q�J����ovR�C�Znm�u��Y�p�����0x/�h�.j�,�3*	��<��ݠ8cڔ���$}����{��aD�e!0�K�_3#ڸZ鎬������$%��kg�ҿ� �,KW�*�	S���{��@-���͸Y֦rVPis��*�!�NrY%T��BPS�)37J*u$)6\��m�,|up�LXS�r��g},�õ��Mn���n���b��1�Jѳa(􆿳�7�pf���ca��H����*N/�p���(�
t�ژq���U�D����bN��ik�&���9�dMbZ鎬�������(���<)G�9� �H�HoLf,0=]^	�&<��)�A�'RW�xAZ"�V�p$��z�q]ެR#G�B�S�[*�$�ᲆ7�l�:Q��Ig`i�ҋX����0�a1i~J��ɩ��-��x�d!��dz��eU��N���\)Ji?N�l�|��].��'���XwM�B�F�ͬ	[�z�IY�/8'�L
�2�Ot�Hb�%�BB$�W%H�˯u�1uXϵ�1��a��B��+��|��].��'���Xw�����犃�8�Qt�z��eU�e��������Dg��y��tqӴ����s��8�M���e���96BD{���p=�Da���Bv�~������]�!�����#e�?���Qz�]�Jg����-c �ЄW:l�mq���)�:;o�������{���_�G���;�Ζ"�љr1c�,�[`�9+��d@���{l�f|����%Hl�(bY,?Z1~�g]�I���B��&���a�%�j@c�rn7Zմ#&<D���l[�!'lBv}�j�-�dnBD{���p�պ����u�Q_�}{KS�)37J*u�v3���?|��(AXAu��,2�����^���@�d�_C�VJ����̕���(��h��1}�����ei�5/U�rQ��3c/��!?V#$~@!<��z��}�צ:�)s�DnV��B*�2���u���d���=A�2�S|���f?��� <9�G��1p�!���j�-�dnBD{���pE�b�.�.ov�~������]�!�����#ee�0��`v�]�Jg����-c �ЄW:l�mq���)�:;o�����p�ǔ|�b��������$�e�7P��T�<��z��}�צ:�)�u����6>�B*�2���u���d���=A�2�S|���f?c%5�H��ڰ݉ �'���ubޣ�mV\�C���osq��|��].��'���Xw�Wl
% ��)ʒ�"��/8'�G~+�3;��\���\ ����@���d}�80�[X�b\g�8>!��J�0N�
���	�Bz���tU`f�g_3#ڸZ鎬�������(���R2�sW��t_-Z��T�\ ��r���(<�u#�ڽFrK���,2�����^���@�K��4��ǯ3�4������_ 	>��M���5^sc�.[K��m�r�������whk�_�בa��@IE�U����S8�����)�d{[���G����"X��[���`m�ڟq��Z1~�g]�I���B�龈4��G	������t4z��w���*#�IQ܋[���,d�܉-`�6�b���n�����띚<�7�6�vg;Je'���Xw^���N�Cp!!v*!��u���d�Ӵ���)�jj���|}�,J�l�/m�	%��>��m������́����H���ɫih��Ѯ��1� Oag�qod�֓��Җe���Z��tveZ�CH��z���8�n��$���Z�"z!��t|Y�f�s\�)8�o�}�� �с�"�,�>E���"5� �S�jn�Ł��}~�oy��E����F��Op�ե[��>Ol{�b�;��1����<����K����ex9f�ٰ�Ř�h�����5	��)��8'����y�]׽Ma(Fj�B��+ H7�ܥ��2�NTګ'6�"z0�L%�B��7y\��<6��$)K�E����F���8�TP��o۩��WM'��9X:i#@���%&p&ĩ+�4��y�'^�"�,�>E��<��z��}���<���_j0*����.1mx���!M`$z�k*�J�y�Pa(􆿳�e�&���6���E��.W�q�1�\�S�)37J*u�,�JL���%d'\�'��FD�ўB�����5	��]�!��5��E0�%����x�f7﹏N�By3��<Z鎬�������(��｀$��G<�K��Q����`y������L}q�
z�.�M�����
L'���Xw�j�7����5@~Ju9gUS��;A���|�+�� VU+I�eC��D>����S������
�):
TTTW�+�@{fT��T�0v��.�/'�����WJHn��z��r9�3]��Y�,��M�P�zL͊�q��b�w�H��{\Jy`w4��#�zL͊�q��!�Vv�P���{ƨ���� w̭G�{Ңn%v�~������]�!��	Ǹ�y85���s#%^�V]��}R�wX�ՖߩJ�9��č�Y���S�)37J*u)T{6T'��OG��_3#ڸZ鎬������E�^��L�����~��|��].��'���Xw��g��[�1��u9j1�f<��z��}�Q2�+�Y�wZ K�Ϋ�v�~������]�!���sC�)��+������!n}y���q���U�8c.K����Ig`i7G#+�ǟ
��|�6|�+�� VU+I��(�@$.>�~�Ι���H(Ť"Of��3f]Ǎc���L7ܼ^GI��'�,����|#^�Vn�^ֻ����XP����w��$C���2c�'z͌4s+�ny�X��{��ܛ�	��|��	(���zL͊�q����#N��RmHX���2c�'z͌4s+�ny��#_��Y~��`�JKݗZ:���'n�^0o�'�=��d&(C�#�7#^�Vn:�}��E5��*��w
j$8c��� 8�2s�. �͌4s+�ny��d�X7Y'ʯv!	��q{�f��a�:&�>��s`�H_�U�A�I����cD���iZ�;`�XHAYIc�V~�Y�T ��7�8��qb�'t����U��R��%�r���c�ż�\�v�[������ڢ��({S���L�Y&��g�đ\ea�G���6(�7QVk��S�)k��'n�^0o���d�p�D��Q�·Τ��ޝsn5d�rfR,)6�h	�q���?˻D?�]���x}���&�����ܴ�&��'n�^0o�X&���5����`Kx���T��<�^0� T2��zL͊�q��e�[,E�Ћ�l�T�Q`��J��k�=[�p���^ֻ����XP���||�?�5�~�!"�-��Wq�;5�s*)F����'n�^0o _xB�I��'�V^[s-�H���A��d�;5B5Y+��
����uK�R��K)�����(�x���T��<�^0�X�I���=�sEټ����6+�y �v��7ir�;��ä����ׁ��m�{%�1%������͌4s+�ny�8b@s�?�D. �6�@Am����;5B5Y+�Ȩ�� "�,|up�LXSP�����q��w{�XW: ���}(8 �����L��F{��O9h_|�9�;�X^��s�`of�i����]���'d��s�KT��s=q�SV.��������=Y��_3L��'9���_�sL�j�赒��_P�� �fb� �1_ӧ��\�Î���Y�ֳ,�Mf���9���q���U���]�G�}N�vʉ!;����K�Q��mm|�[B�����'���Xw�P>a�.����'�#&�3��3���$�],�i=O��s�j���dDqS�,֍�Sx�lޞ�-�`��8�4���[!o��Ļ���p�ʅ<#"	7�B�>�p�:�{K��q{���1H����Ig`iZ鎬������=X�~���X%���xT����^-�����G���;���W�v�T�
nː����[B�����'���Xw�P>a�.����'�#&�3��3�_��PN������;Q�U	t�ޤ�
�_�[B�����'���Xw�P>a�.����'�#&�3��3�~�̳o�����;��K�Q+���)Z�O��=Y��_3L��'9���_�sL�j�赒�����7��}���D]򤰷������K�Q�c��Ҏ��=Y��_3L��'9���_�sL�j�赒�^ŇI���O;�2��~=,������#Tж��SF���v�Sx�lޞ�-�`��8�4���[!o��Ļ���p�SBc�8��
���;򤰷������K�Q����-/�Sx�lޞ�-�`��8�4���[!o��Ļ���pD�?��#�H��õp򤰷������K�Q�{�<��G��=Y��_3L��'9���_�sL�j�赒�����7��ǡ�����sz����Pq�ҷ���� ��g8���D|-o�Z��beNY�_Q路��K�b|[Sx�lޞ�ό���.���K�Q�f�3�Ұ5ϝQ��������B�['���Xwa'�<� \�_Q路�/8��A0�1��P�߭Z鎬����D^Rm�	�C�<��F���Z�-���&Tʥ-�
�W^��P�F�M��n�b0���=Y��_�0z�cULOE��
��x��±eKr�V�fR�1屖ʨg��U-�e9��K哧-�
�W^�@���°�E���V'/Sx�lޞ��rs�i��H���G��x�#���FU:�\2�O����	a(􆿳���t�$���JL���Z'�A�җ�*Mf���9��Y�{'%sgeߪ�{���b�QOu��
Q��x�'r����MM
��,=�|.�Tӏp%����l�_��^�ȥMf���9��Y�{'%sgeߪ�{���b�QOPǨ�o*� 7�v�ԯ�o��f��)�`E5U���c@���G��Sx�lޞ��rs�i�J�{jo��,|up�LXS�O����	a(􆿳�>d�ˤ$T��@$˺/t��꫕qŧo��K�O��C�V�j"���C�t%>^��?�y��hL5ӥ�����B�\K+����!� �,J3�1I�؊�"�D
e���4��=�!ߝ��X�!� � _����J���_P����b����";�S���o�>�5�ﻋ-���C�M��N��B�)��x�ϝQ����\Ef�>�Q3U�eT(�q���U�)}zu��`����׫�Cc�kbi��G��[�֔(
ݪ	� f8�p!!kU�7�X�3�ﻋ-���C�M��N��qg2�K?\�ߦ�����?���*gaB�d�٣��c�A�L'w�d�b��X�Q��[�'r����MM
��,=�����x�S=��O7H$�DZ� C�C�.�.�:�L�
�+f ;+/���['���1�]�!��	Ǹ�y85��־���
��-���Zx��[�Fc�k��`y���pzl��a�r6����b@�U(����=Y��_�0z�cUL�?d�)SһN�ʁ������BT�^���8�B����`m��8�C��lŨ����R�f7�[�}��|:��T�]�	�_t����?�f�����}��Y!��]�!�������DTfF����%2B�܎���U�������K�Q�A�qL2�cP/���[}��=Y��_@D���uL�ɱ=��C�o�u�/@&W�3!Pc�1�QQp0��J�˚�Jz�0���je�Vm@�Ɇ�hq��P$��j�t��@a+����61��7a	�����Y�
��LG��&�'�3�$ �#^�Vn[)�ٽ�f퀔�������sr���0G3����T��i7��+:+, ��ɧ���7�)a���%}D������h�br���lpda���\��6m��B��${��?�J�Z��]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gV��Vv;�Oe�d�#���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���))~�� ��-[�v:v�o���+����7X��U�?	r���/t�u�9�GKP�2�����Vcv�iL�D�"�
����Z�q�PO4�:_b�b2�����Vc2�����VcAQ@;�(V����	�S�J9!�-� e7P!*��_ӧ��\�]�~���S2aw��N����b�O}��XHg�}�3*±�)c�>�ӼM�6ޱ�|x"$�.�;�H���o�QuU����t�&k��@�&��}s	=Q+�����3c/��!���M�I��s��I� �/r�[�DZܤ�j���ǈݻ<6}�~m\��s��IȰӥ���C�;�H���o��և�GIt�&k��@��u8ۯ$gI�3]�۞h�G��e]�ڭs,��f��=Я���)ͼ	=Q+�����3c/��!Z��19� -J,�ɢ ���7��Ѷ�DZܤ�j���ǈݻ�p�7$m8-J,�ɢ П�bWVzH캧xӍ.�ya0���U,�E{�n�����ٹɵt�5W�#�v�������ƍ�M��7ì�����$�'DV���b�z'hۉ)<Y��=p�
9�GKP�2�����Vc2�����Vcl��w&� 	���#�|"ap�� s;���*5���(ZH4~��2�����Vc2�����Vc.�
͹U��|"�I\�D��y��w�Ϛ06d��-�����R���Mصd������h�1����ԡ���كs_����fB_D��qh�;P��Te L�J��wfl= |P���Ϛ06d��-?^�é�;��	� B�\�B+]L���2�����Vc2�����Vcƞ���tL���f��#�hr���2�����Vc2�����VcSd�*-}Q�g�}00
W�Vc�sNL3�ͧ윎|\#��Z贯x�#���FU:�\2ij.!@J%A�M뵨�I6�j4̗��W;��"r뾃	��s�G��,	��=7)-/M�5i$ۇ��;"�1���dUl��3c��)��HS�Q��[���$ܦ��%��ό�;�LȫԷ�/�"�Y�%u��h�}l��F�����ٕ�����dc�@z�ׅ�ؘ��N�g�c�`Ѩ�f?�R��u#��y;��"5����z��c� ��*��؁P�y�����S�T��=7�}|��	�/̥@X�4���'|b<���1��X��WG ��U�L�{k	�#�O�o[v<�F����O�%U���c@��`Xg?�g��z7M�D. �6�@Am����^�V]��}u*w�A�X�H�->t��w#o�]�ʄ�"�G~4��9�ͤ3�8���~կ�@/��r ��JR��W�xU���c@��`Xg?�)�$z
�*|@���°�E���V'/��.�[ ٓ���>q_W ���t��������*=���$G.
�=θ�=7�}|��	��a-6�Da/8��A0�T^���!4;�gˬ3U���c@��`Xg?��i����w׏�����MJ�1���۪	�}a�]�w%�oφ��<�6��\���BP&��T`��J�^E 6acsO�`�;MV\��@�n���c�SV^�V]��}%鯅�W'9hha6S���";�S��_չ�ŉ�T`��J�^^�F�_	*�`�1v�-�/{�3C����^=�����l�1C��(�H/�I���΁�4���p�ɟ�V@�]V�g�}00
�-�=5>B�úkE�Q'�)r�E�9C�����dcT��NB�D�u�<�2�Ҧ1���Z�וzj7i�j�L�4�� �{1���r2� N��r*7O��4'أͽgF"?���b�QO��:F�X?o���wu6��V(�z%aVW��
��{Ba�nl��+ѝ��WT7���=�~���i�xM� t��φ��<�6�Ps_*�GqW�w��fDT�<bi�[zB�L�[���8di�?�{Zk_.oʛ~��"�����n���wH�-��V�F�P�_�^���\�}/8��A0���:_� ����O�����S�V��,\ަ�It}�0�.�,U��G8���z�r{]i�X;p`����b�QOh�{V/0_�=2�N�{u!��}.��}@",|up�LXS�c�@9V��S5A͍3��d�)Î��C<봯x�#���s�3��o��~�;����ɝ\�!2A4��y�'^�.Y΄�l�jyd��- ]�//� �c���,.Y΄�l�j_:�VIͽ�|*�>-t>�e%�2��l�@jen�-���<8(�?Q�=7����U�p�6j�"Hs!�pL_��{Zk_.o��AZT	..�?�ۢ�=e��6�Յ����hM��0�d(_\�^?'qKy���\N}zp�jN�W%m�������j_P b�5��Eq�`1�
�8jYj'�EI�[K�f�
�`�*%0����W�������9{�?���\@��u���?�5CJ�ݨg4$`�^WZB�����ɧ�+�d�_�t[ⱸ�ND[M:b������2F��uP����.(�o�Z���h�WV�#a�H���w�@üߦ������-�z@/8��A0�@zS�WV��	��y���rk���&�e���Fc����7���z7�|�|<)����j��2��~���X�<H2�W�(F����}��� ?�d���&�D�;E���<�����&H)����g�0�u��a�֧�I��3��a�����x��L��M��liJ�9J?�"5����6ջ�[�^�T`��J�^��,����rw�&�z<a��N� φ��<�6�t����˴�|���d� ������TU���c@��^Q��m�!Όg&W�w��fD7BP�m(�*��T=s ¾@\�j�'�Hm��1yu��mDrv9��}�c�uP����.(ʪy�� /���`�n��U%aWp��.�替��+���<j�2ʧ6�0�U��{L���D5�p��.�	�ZMC3�?�AO�]�����>L�k��cIEw�S����?�&����]�w9"x�g�Hz�Ó�[���2�����Vc2�����Vc��Y7���$���K :<��ޫ��8���N�1�� ��2�����Vc2�����Vcbc�~U[f8�p!!k�ܒ��+Z�T`��J�^E 6acs���@�_�c�x��±eKr�V�fR�1屖��i����4�fg��e��ł!ڕ
��+�^�dQ�3L� n2ϒ�ȃ���A�ڈyܤ�܎~��$��/��^�<de���k	��Ո��sZ<�����W�}�:�Q%�h5�'����'�2�����,�>) n2ϒ�ȃ���A���@F>.���*^������CU߈!��A���ڴ�>��XO��C��SkXKWT�����	��Ĳ��\�uB�3DO�9�?��3LO{���)�u��ݵdw3{����kGQ�����_����7��EEw�S��EC��Us�_��s�֙f����hڿ�����F�ߦ�����E2�4� n2ϒ�ȃ���A��{��(:/�b�&�q��p�Lu��z1h��ʠU�n��,3q�$���j�/A=�8#�H��7Q�lՖ�|���d� RQR7�f&���˓#���2�8�Ǯ� ��SD�-�e��0�UҸk�2�Ż�&ǥ��a���F߸��S�Ȍ��"+VqS?�d���&��9��^K��7�H�8i�H�玨���8$���¸_�p�u�aӕ�:1�	�k	�8$���~��"����(t�	H�޹q��7<�|ޒ�i��̋8��syu��mDrv�H���`?�d���&�D�;E��Aq�:�5�`_�ʵ߹�)���1h��ʠU�E�?�j�B� ��~��;�9S���WH�b�y?3NϜx	0X��f*�a�	�+4D@5b��-��m/�J���I��nF���	+E�5f���%�ç�˓#���2�8�Ǯ� J���-�fB�^�4,+��77�4ŹJ�1���۪	�}a4����@[�_zβrꢯ�wv��\�j��fxŪ5ex:���t�eu,00}K'���P���]��CA)��[�uJ8������CO�$N�F�J�O��")�/K���i��vp�Of�,�8�2	� �%y�7��0Ba�N�-�%��1gkQ��@Ő��t 	�J��Uo;xw��i�6YF�1����GL�!����%���V�/��.���oE��)L@�v?�[��\n@�>�~������b�d}�.w.cҭ=+�~��"����(t�	H�޹q��}����M��̋8��syu��mDrv�<�2�Ҧ1���Z�וzj7i�j�@���-�qx�'|�9��x~l��Uh����L8�C�	R�x�������ՙ�.�h͉��7,F��[WL��g8!�|!��[�N�g�c�`�zc՝Rq�	�!٢�,|up�LXS�O����	a(􆿳���[� �G	B�^�4,+�����l�TI+a����R�1屖ʨg��U-�e����k�l�[b%Ɨ�������ܻK;��I��=�sEټ�*��T������z���nF���	+E�5f���%���5ߧE4��\�ܢ��,	սL��$����,�ǰ��[2���PZ~���6�틳es!FּQ*�:1�7!p�!��I\+�a�/O]]u����;��9C����#;�ec��Uioέ���'*$�T�n��
��4�)�� G�/�z�)�_��s�֙f����hڿ�����F�ߦ�����E2�4� n2ϒ�ȃ���A��{��(:/�b�&�q��p�Lu��z1h��ʠU�n��,3q�$���j�/A=�8#�H��71ri���ђ{)8A�^�V]��}�dh_��tCdN�<@Iv����-�T�8��e�[b%Ɨ�������ܻK;��I��=�sEټ�*��T������z��|��*��'|�9��x�Îa;�`ђ{)8A�^�V]��}u*w�Arw�&�z<a��N� φ��<�6�Ps_*�GqW�w��fD!��I\+�a�/O]]u����;�7�u�l���V�{��\|��EaV�5�j��K�����6����ɣ��؅)�{�/���`�n��U%aWp��.�替��+���<j�2ʧ6�0�+$OF>�X����Y ����-	��ȥ��%��VB���/ r�F��	V�����|�%����_�=�4wW'/���d}��[�ƭM��P���?2�����Vc2�����Vc2�����Vc��Y7�q��$]�W��	]�	)�(#�� !�hr���2�����Vc2�����Vc2�����VcAQ@;�(V�x��p���%�$�zr���įէ3[�?�����l����4�n���xǊ���PU�p�lJo:>M�A;��h��(Z+�<Vo�eo*�ڰ3�%c��ɣ����x����>�M��K�2��Z^��:�S��m�\��jT�):1�#��йGB�����*rcm� ��>ar��{�&���R��K)��u��p����K�)�PMI������NϜ�cb0��w?�h��(Z+�<Vo�eoB���"�zђ{)8A���,�am�^
L�PX~��yy���H��+2Ph��(Z+�<Vo�eoB���"�zT��<�Ux���T��<�^0��b�;���Q��m�f ;+/���]ڨ����s�<�i��N}H����	K$�ْl��]�B}Ю�0�`m��';��?2^�9<o�nïi��n�5�F�^hq��:�����+�nt�x��h���X �V^[s-�H�	�dV�Fm�#nS#y����m�zЦ�+;4#`[�=I4�����	T�|�lSԃ�N�y�@~�MԲ���d��#��R6�.�ap7�L}��GN�`��B�0w�>���4w�g�P_���7�gI����I�}jZjx��7~���Ho�d�	r������oE��cFl����h4c�H��Y�5}٨5�X��o=��i�h"r����SX�c�,�[`�Oʕ3>x����`4�E%h���R�ނ6�l�yŶ��띚<�7�B"�u�������D�� >r�Z	��R��	π2�����Vc2�����Vc2�����Vc��Y7�z�p���w����	��-�d{��%�|p�EN�1�� ��2�����Vc2�����Vc2�����Vc��G�ZB��uB=+��A��寗Z��/g)w������?�7r���g��%�fQ6�F�����ٕ����1 �u�.�a�	�+4D@���^xc[_3�mE�_se�!���@p)�!,�!�R��q4ً�?�(�p���� L7�i��6ð��T��/�ciJ����	a��=7�}|��	��a-6�Da�A�qL2�cݽf�i����Rh �rw�&�z<aSm�6��`4�04�jf�5ߧE4��Fi��|�3;c�<Aj�X���W}sû3E��|�}VꌗjO�����v���f��*c>��3DdZ0o�vʽ'��G"����6�M^>�|�uI\L'�+;�^�~�祠4��r���u#��y;��"5�����Bl(�Y��\Ef�>�8��W�%	�#�O��)�	��r���|-�se������D�{�I`�	-�_3�mE�_s�rp� �1x�it���w~��,�F�,����1��X��WG ���zt��[��t9��\�w�xo�A�\�G���o����Ӫ�/8��A0�Pع���a�	�+4D@��~JFN�wOm���	�#�O�o}����ĳ�e��@ai^w&����|-�se�Pع���a�	�+4D@��~JFN�����J�x�Ǖ[�Ps�w�xo�AB�R���>_�;�z�3���L=l�(��|���h�x#�L_�(D{ͬ�y�4����Pb�)b}�FL~΄gO�3f��*�����R����b