��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-~09h�i�Nq�{5��]�0�lK'���Xw����Q4f����om2�YQ}��1\���^�9:�M��z�}�I@�;摼ڃN\��~�����]��i�i�n/�NE��l�JHn��z��[�Q-�͌4s+�ny����@���_�G��G;5B5Y+�Ȩ�� "�Q��wjw�K؞FMN�*�])������u���B��C�QU��}<o�Y�d�*�K�
���A�F�7���3�GXS����E@��~���($�J.���
�=W�֯�^��N�&��?�2�1p���}������]�0�lK'���Xw��_
�u�m�\��q�Z˻r����4��a�&�������N�N���aC�h�>W����Q�\DR]R�x!���2͖梡���h`�fx*���-the���ʝyzL͊�q��5�?����F�U8�3���lHc�,�u�:��ܣ|4�/��ӝ�9��,V z�J��x�]Ҙp��0c|=}�? ��i�+���9�)bv'.8��>oUa/�OZ�5�p�������m�X��Y�$���e��y~}�;h>xQ)JC�4];ˍH�ƽ��s�I2�}1R$Z�#�u�q8�6K��uIm1��y��/e��^p@f�Ԡn�gg�L�@�1��ꓩ�l;��!I/�������A��1��+�W��J�ݨg4$ _o���6cMH%�]�<o�nïi�;5B5Y+�T�����NF@��u�'�3�$ �#^�Vn�;ۂ��IÙ=�H���0�EѠzM8%�Y~��`�J=�C��a���\�vūx`��:���Ϥk�;��|B}ø��y�w8#�RC�G�G~��6��m:y+������pW�F��F�zL͊�q���}o��E��~��0�#Z��pޒ��w
����2$6�sI=�I�Q��u��m�dR���8R���|��J$���I����`��Z��@|.�dkc�;ۂ��IÙ=�H �:`֯z;�=����ҶؤƂ��l�'����ںV�^�Ez@y����݂; ,@�� W�h�)cGO9��< ���!���Lʚ����9X�_K���1ƚ,�0���^ֻ����XP���ĵ;UQF����5^���L���UN螗T�2�K��G����Ǚ�*�������:�A?Љ'�-��<v5b75�H"�wZ�pC��)Va.E�}�.�C2�>d�ܡ��5��8�t��\�v�x��L�B��:�ʟ�����R�fPذaf��pD�Т��?�(j�"�A�#�ﷵ�;�|�:=�V�	s�A5X9:)�׽�P�d�����y�:�B�t�LǜI��Ω��n�[��Ig`iZ鎬�������(�����>9UW?8�����m��6��Ԋ����[,�'��j���^N��Th-h�x��pc �Y��bp;�ঔ^ֻ����XP����Ql�Z,΁��5^��t����
�E[DN�����0a�b��:�m�Y���K$Ÿ&Ot]�ZxE�IM9�����S���	����&�6~ [�Wxr��U�KT��}�����FQ�03�^	�[0
��{r�X��B�W!88�L�� �E�<k%���d����l��Q �!޶9k:����2��O�����qθ����;�� X��v4��/t0P_f�$Y��X�W�F��F�zL͊�q��G�D�� �~��0�#Zu��^��.���o���
��/j�~�*�.ie��-�	�hZ63S�݃O�hf>Ŋ Ύ=}j��֢8�٪3����?;5B5Y+� �i7�sp>}�-L��-�MR��[m�>���$�_o�EO�Htv' ��E�8h�4d�>�/���8"'�y��59x+�	����b��X���n�O*%�����Ϙ�M�o�^���z�0�>��	�Υ��9�dMbZ鎬�������:�!֧m�}`s�4��<�K���>������<E�Ԓ�WM�%�+��gӋ-�;ڨ5W��_K��8k>6s����]�!��	Ǹ�y85�R̺�?})u�%N����`y�������g�EH�a���sbbj�i0�i�G��'(�R��G�
~H�>������<E�Ԓ�WM�%�+��g.�p�c�#�/yص�3n�l��\A$r@IE�U��|P�����@�Ut���F���j�_������ZB!g��nB�nrm؊(�o�@~z����v�h����~��4�Uك�["�x�;}�z�5\͘y'��BS�s�Y��A�^<�ҋ!����8f%�8k>6s����]�!��	Ǹ�y85��3}�@�7	s�A5X�g��U-�eRAѭ�����Ȧ����:��
K]}����^<�ҋ!t�}3k30�|��].��'���Xw�j�7��ޒ������JoEѰғ8���/����mm�<%l}����Z1~�g]�~����0_���>���̈�1�WC��nk����Q�Ar+A=n��K�//�����c�9�:&�ߦ�龔�Π��č�Y���S�)37J*u�v3���?u�e�+����nU��\�x�/8'�a;h��ά��9�p���ٜ�U�n~q_3#ڸZ鎬�����r44���ڶ�|ceJ�z��eU�e�����T�2���%,J�l�/]��-5L�8`�#�I:)�%����7����č�Y���S�)37J*u�v3���?8cR�F�㯆ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,�����Vt�%����"��#����V�a�QtDo~e۞h�G��w�O�r�e�!n}y���q���U�F��Fy�. ���ѡ�e�LZ\^�e���Eы�`�M7Э���j�ҹ���9���ϸ�Q�E�"�D<��ͻ�U�ES}�T����3c/��!�{m�
�<��z��}�צ:�)��H'�񽂳B*�2���u���d���=A�2�S|���f?��� <��U�-�R�so�	�C��ypj�p]��9�p���e'��ǩ����l�u+�v�~������]�!�����#e���J�l�]�Jg����-c �ЄW:l�mq���)�:;o�����G�̥}�ߘ����N��t.r�������� mc�,�[`�O?n���{l�f|����%Hl�����X��Z1~�g]�I���B��&���a�%�j@c�rn7Zմ#&9�� :ܝ}���D]g^�*����)�%��4_�;��	�ya0���Uu�Q_�}{KS�)37J*u�v3���?�I_�=0<��,2�����^���@�d�_C�VJ����̕���(��h��f�<�K6���x��B����.J��h�D��0.�Q;�m���|��].��'���XwSn����P>ea���||��/8'�G~+�3;��\���\)�K��b����(�u�b�)���8�V������ͻ�U�.YUr�k��7P��T�<��z��}�צ:�)e�>��E۳B*�2���u���d���=A�2�S|���f?NԆ��-�ê�%�S��!���A���ՖC�͓Wԙ�"�F�%d������hڏ<K����>�Cb�|��].��'���Xwd�n]N�h��7?����Wǖg3ȓ8���/�G}�tL�x�N=�0��]�Jg����-c �ЄW:qBbr�a��\�"ߗt� ��wg|,���%�̈́T�٥��T�%����@'��o�/�ʹu�P^��*N/�p���6�vg;Je'���Xwd�n]N�h��7?����Wǖg3ȓ8���/�G}�tL�x,-6�41�e�LZ\^ �@'�ZX8�5}7���_UVp
MMo�����!Au�UO>���)E'��o�/�r�3P���WT�j
�I��w��,Y�?A�3����a;�/8'�L
�2�Ot�ky����R� -�*3fN&����6F��ŜgTKfVutְ0�]F$�J�q㧵�0��]Қ�Jp3H�Q���,���r�R�k&���#�{�0;�}�f���R�\DR]R�x4�mm��Ix���� �~��Z2��u�>��{=��[^T�d&(C�#�7#^�Vn�^ֻ���(_�<��+�nt�x��W�F��F�N��B�)Y�l���n�2�y�� �sq{�f��a��ͣx�`&}�K�
�4l�G�pޚY�i}%_3#ڸZ鎬�������(�����CcO^Z}��"X��[�`�L�i�GV��y�&_3#ڸZ鎬������e��9���b\��!n}y���q���U����c)0k"�Ι�y�Ң�{l�f|�ό���.�{�:���g��č�Y���S�)37J*u)T{6T'����f����|��].��'���Xw＼.o�Þ�7P��T�<��z��}�Q2�+�Y���R"@ПWT�j
�I��w��,���|HH9M\��e���S������
��x���ӄ�bİ�����ap�]��5��f��&��$�B�I:׷�F׫�J��q{�f��aƨ:bN�t�ɹd�'��"������JI��'��'�3�$ �#^�Vn�^ֻ����XP���8TJ�����[T�)��������JI��'�@���U@���:��F���V!���IÙ=�Hٍ���]c�PƐt
�2c�'z�㴬]|~TdZ0o�v�3�Dc�`��rj���9I��'������R�ê�C����\�vūx`��:��5����`K�b֨#u��!7��5;5B5Y+�T�����N1�*_��ha�G���6(�~)x4�;ۂ��IÙ=�H�\�'���=�k2B]p��	�/T�F���}�� JHn��z�IC��]/?.i�����q�f�7���n��b=�kM4v/�?��_JhI��'�f/Dq�)�0�y~M d�8q{�f��a��pP�o��Ik�v ���כ�?n	�����>]��|��~�Ӆ"�5͌4s+�ny��d�X7Y?#OF��KݗZ:���'n�^0oLAfʶ�Ա��ۖ�lhllEۀ>7�͌4s+�nyL�m�_�����K���nU;"�~[��\�vūx`��:��5����`K�0�Dʒ��d>v��,uYL��ٿ�JHn��z���G7��͌4s+�nyL�m�_�0���2�W�ub���<p�T=���e��IÙ=�H�\�'���=�k2B]p�^ǙPn`B]z(,ߔ^ֻ����XP������DK=󕏜9����F.�!˯﹈�iq{�f��a��{oS���%�a�e�ٔ�"_�ct�:��RE�$<���GzL͊�q���`��#)y�I��'�V!�"M�Ϭ���!I�;5B5Y+��q	k���A�+kG��Y�9��'EoU��՗7r4��c�����\�v�)��+�}�͌4s+�nyL�m�_��"�m���r�;ۂ��IÙ=�H�, �dh��X+)%`d�Y�Y���҇;-;*�7���|���\j�<lG�"*���.��F.�!���LI�.�͌4s+�ny�8vZ����_�G��Gq{�f��a��{oS�n�1:`R<^���1���3���!�͌4s+�ny� o�������Ɲ&�Mf���9��Y�{'%sgeߪ�{ޒ������JoEѰ�MM
��,=F��Z�ؕ��������Wz�p���w��Z�-��ݾNt�Y/�n�*���}��U��Ř�=Y��_3L��'9s��j�ŉ�h�9:De�;.��{C������������6/�
�Nyy;%a=�'�
�h1��	���s=q�SV.��������=Y��_3L��'9���_�sL�j�赒��_P�� �fb� �1_ӧ��\�Î���Y�ֳ,�Mf���9���q���U���]�G�}N�vʉ!;����K�Q��mm|�[B�����'���Xw�P>a�.����'�#&�3��3���$�],ߑm�������K�QY/����[B�����'���Xw�P>a�.����'�#&�3��3�-��y��hi=O��s��#%��$�z��e�K���d�٣���-��� ��d�_C�V��pµ�Ս��������K+I�\z�f�a��c�������7P��T��]�!���äs_���l�mq��L��T��>��Nv|��U+�ei�N�iP+����
�_�[B�����'���Xw�P>a�.����'�#&�3��3�~�̳o�����;��K�Q+���)Z�O��=Y��_3L��'9���_�sL�j�赒�����7��}���D]�A���l_-B�g��^�z��e�K���d�٣���-��� ��d�_C�V��pµ�Ս������5�u��z�f�a�Ո}�nNg��7P��T��]�!���äs_���l�mq��L��T��>��Nv|��U+�����N�iP+��w��n��y[B�����'���Xw�P>a�.����'�#&�3��3���<�4������;Q�U	t��\�T~�SMf���9���q���U�?�����"2�#�?�< TL�MK}�V�h�;����;Y�hg�N��M���5^s��Z�-��ݾNt�Yӑ!�;�?��R��V�
�]�$��'���Xwa'�<� \�_Q路��t���(�xw����$�Z鎬����Y�V��#q�e�1H�z��T^���w����$�Z鎬����Y�V��#q�e�1H�z��Q��ٹ~��ր[��d�٣��20X��"8�kѶ���� ۗ;` �ܑ��݆Sx�lޞ�ό���.���K�Q
�M�j�����[s��� �`V9C�]�!���o��w���tt٭zꡍ��>��{�50�Vr�t������j��9����G��s��d�٣��c�A�L'uab#oLpk��Ǌ"�G\O�E朦�T�\ ��퍥6��n�\l쎭U(����=Y��_�0z�cUL�ȘB�k6~.jʳ�R�1屖ʨg��U-�e9��K哧�	�_t����?�f�����}��Y!��]�!���o��w���e�7-�o�� ��M�����%Pq�^�)}���/�|_�������)�'A�-�Sx�lޞ��rs�i��ߖ� ���y�:�B�)u�%N�ߌNu�5=��<AUy�Ţu!�y�2�z�S�Lw���7�J����=Y��_�0z�cUL=�[�A��������p^�V]��}%鯅����?������p�'w�I��'�1P~9V]�)}���/�4]d���z�'r�_�(pSx�lޞ��rs�i��ߖ� ���y�:�B�)u�%N�ߌNu�5=��a'�<� \h$p6��0Y d��W&�]�ר�]�!���o��w����KxC������H���Q�	wM�M�����G��[�֔~u!�3Vt�>�z��^)+��ﻋ-�����S8�<������K@�>��C�4�g��U-�e9��K哧~u!�3Vt�s��1^~��O�$+��ﻋ-�����S8�<������K.?��.7�,0=]^	�&QR�u9�����K�Q�&�������_S1����9(�Hv�������Y�{'%sgeߪ�{�LEh��� �Ne�^�V]��}%鯅�pzl��a��m�6zi�����9�tI$U��K{~��usZ鎬����Y�V��#q��U�^���nRdd��"iNQi��]�!���1����m�6/z��jv�]��a����g�o	�d�)�q���U�pzl��a��m�6zi�T^����4D���t�2B}G�J�ό���.���K�Q�&������(N\�(��`���ݐﻋ-���C�M��N�۔�Zr�X�ȀY;2deM�|�2��� �?g�Θ�Q2�+�Y������bp'oC�X(_��89|����gV�hx�:@��]�!���1����m�6/z����s\���o�e
���d�٣�����6>��~u!�3Vt(t-�D��ht��g��8���O�'���Xwa'�<� \�j����flR�����i��P
Z鎬����D^Rm�	ʿf��_��7�
r�l��Z�-��ݾNt�Y���l�f�`�`Ƅ.�$E�����'���Xwa'�<� \Nu�֧���k]m��Mf���9��Y�{'%sgeߪ�{WW<����,0=]^	�&QR�u9�����K�Q#t�,��r��WdM4@�.'���jJ��]�!��	Ǹ�y85����S)ÿ�M*����9�U.��͢�����S��(�M�U��V��٪����mj�pzl��aꬫ�;�Ӏ׬�����D��~��n�'���Xw�%�fĀ>�[<cP~�t�%��ͺ#�[m�r��ٶ�`fP�?���&<�(v��2�uB=+��A��寔ݾNt�Y�{�W~�_3�mE�_s���R�AZ鎬��������}������$h��qa]�݊3�;|q f�yv<�1���\�۟�-?�d���&����{ԕ�/�����jt���@
�ѻ��`���+=����7�>D�c�lQ��� ����7끍J�[T�)��b�����6��`�n��U�z��pU6�M�S��2�{��΂��1\�����s�[h}�k8�5�>�yKYQs��[�|�F��˱4���[�jDG|��o"� ���I��Q�yt�G�^����]S�WI�;�_�	�t쩖NUD60L����L�Y&#t����n�~����p��l�n�Zlmך҉ݨ&@)�F� ��FZ���;D8���:��M�S�ᳰ��X�z���t���Xo޲G�����$7x�c >��}f]���]�w9"x�g�Hz���MN����!I/�������A��1��+�W�Ń�I��-Nd`*3�'�&�2�����Vc2�����Vc��Y7�z�p���w�nrm؊(�p��Aby�2�����Vc2�����Vc���1� -N&ݨ)�����a��	{��#-�	=��>QH[[����q�f��6&1�1�<Y�W�q]=`爼#��8h� 1�����f�c��k�-����B���f�;�>)�(���Yr�r��`�^�qFQXI�DZܤ�jh"r��RǷe�b��1j�L�uVBM�d��_��;�H���o��l�u+��[��U�D��sMO�2�h7�a��c�,�[`�Qb��~���y���������DZܤ�j<�`�hE�c,W� K91j�L�uVB��=��|S���I�&�`��\��K��A!�?2���L�b3N��wm��5�;�H���oՖ�zA!�?2���L�b3N�B�����f�;�>)�� �4"���B�V9��~(j2�����Vc2�����Vc2�����Vc�m7���e�*��w
j$��) �Xy��|�h�E9�GKP�2�����Vc2�����Vc�C�z��/|R-��]_:�A�����q�J�m>�Ф=O��
2?a)��R�����OwAg1,�!�q�J�m>ձ`��NH��l�����dB�;n��
v�Ϛ06d��-+}�#f�!��3�xʣ^�*�ǒړ��Q .�L�m�����*�ϖ�	n�h���� 1�=��:wB�;E��qb�2kl�,�;ڒ�!_m���_A���\�b^
2?a)��z��|B��yk�9��^�كs_����fB_D��?#OF���}Vr	��9�GKP�2�����Vc2�����Vc2�����VcREBR�hHr!޶9k:�������M����O�b�`q�M��9�GKP�2�����Vc2�����Vc2�����Vc>�P��^ez��X}@��M�T��ےOyTg��q)�Č7O�-�� )w`V�;��Qz�#g�k��m��uJ"xO��H{��B.��(lD��&Y��V�^<�ҋ!�<�o�2JC�=�&Akgc`��g���;�%�L
6�,��V�F�P�_�^���\�}+���Ã�*j�xXaZ N��r*�?�I���6\�4�@���(�?<-M�O��~�Ѩ�f?�R�����bP��a�	�+4D@���'9tT4]d���z�'r�_�(p��-x�<�cFݡ/��x����u���oVl�(�!�G}��z��9;�B�|���qbsZ��"�)�{�°!�?����S�)V��B�1%�x �N�t&����1〈)�����d��-��!rϚ����5�P3 C��Pع���a�	�+4D@���'9tT4]d���z�'r�_�(p��ӎ��������Ս*�(f�Kp�-a�D͢fU�9�׏�����MFi��|��wØ�ߜ���,�ǰH7"LTftYD3���L�6ߟH��Ǵ�ԏ'dNT9�H+�C@�Wu�t�Ru�A^Hu_�_�뱬�WV�#a��mJd��?�7r���g��"����0h�5e��`'��<��Ȝx�� BN1l�n
V~$�~j%R��W ���t�-M�O��~�n
s�] �ۆiq�L�ۗ]6�Co4��{Gyn��5����`K�/�����������1�G ?�Ia�fa(􆿳�ܠ��r����s ��,�Y��?�/����s@L�Zao�o����Q�?t�R_�f�Hى��_�
k\�^�sW�w��fD���򫒡�7$�_:Tf�S��6KW ���t�������R�����OE�V|{�@/��r �f4%�!I�y�!��G_	���`Xg?�v[S�d�� �����CO|2�@#k�˟ܒ�o|k�Lb�5ߧE4��\�ܢ��,	սL��$�c���1�ā���z��.��hL? ���U��W7���*����KCg�:�X���o�u�/�G'g�r&������h$p6�CPN'Ŷ��eM�k	�xw�<2%�{��(:/�b�&�q��7x:�����HŹn�M�#�P#^�3�� �fU�}{�h��d��-��!rϚ����T^����H��	W��N�g�c�`�N�����P5�E���E���V'/��ӎ�ۆiq�L���o�/��rG�{��6�y��_#O�/�0׏�����MJ�1���۪	�}a4����xZ@4�׻xO��H{��������{�i� �uC�f�hV��{V�
���{��*{8N��ǆ�K>��/�+�riJ������qθvZ���t�S[�r��@;}�ӑy87�F~��o�u�/�g'$�F�c� -� ��+�����p.��=�A���tMOG�WKj�G��U$�yu�n�D-����p�m~|�֙2{.,��V����:q��n���XmQ3��Tgʱ=�+��c���W���M�;䌚"HG�`�hE\[���H~���-O ��.��G8�H"�I�<�,�+�u���$�n�sȸ�"rR�"nt�s0���a|&�Yr�lc7Bo��Tzj��v��ܑ����V��WP�����m{IޡM�%�|yU��������5����`K�WF��0g��z|5��z	q@��57�1ʾ�!�����@�)�I��F|>��iBM������D-'��7���uD�	|_�������)�'A�-���P�ţ��${�p��XFf��L�'Ķg6�Å���E���ȶ��ՙ��x(�[.��T��?�IdR<3;���#ְ$t���b�l�1C��(�p�m~|�֦*�V$ ��5��4�{Aj�X���G-���6��1B�:ͫ�C��MZ�w�R�H���|
D鞪�%o���w�a��D ML:�h��7?���?eY��5�g��U-�e>� {�}���my$�N���Uە��g?	��oW����
�/|R-��]�C2%�{�� N��r*�i��"u��/|R-��]��A�1Wk}�aá�����-��ol2���a�H��	W��N�g�c�`T�+rJ}?I|`�ht��32O!j����7��|�K�Mv!���x�6/�%���v�i�a����w��ΊB>���<���Hn
V~$2�t�N��/ѿ�����Q�9_*p4�-�C��7u#md��X+-U�9sI�ߋ�\��O��V���1��X��WG ��T�+rJ}?I|`�ht��32O!j����7��|�K�r`r��|`�ht��32O!j����y��m�0rw�&�z<a�4�ڈt׏�����MJ�1���۪	�}a4����0�v��4�����lG�_�.p����P�f ��ME)��ƽ��Ү����,j�W�q�l����K��֍�`n�Pղ�ΥT�t�R��9�u�1It�� ���F.�!�b!>��]H�2?k�v��ΥT�t�R��9�u�1It�� ���F.�!ˆ;��(dU�m��D��*ڡf��m[CMO��c@�Wu�tu,�p��'�'VV%�L_��s�֙��#��j��9���ʨ��N,���K�x���Q�;�hE�ǐŭ%��v��M�߾ol���'|F�rs�(�̴Y�{'%s�6F���y����z��`�"�m���rYj���ط^��Ǌ"�x���|���3U(�{Hl���!#���.�h��&r��rs�(�̴Y�{'%s�Ǹ2����y�:�B���~8���ct�:��RE�����|77*.��]F�j��9��疅(������l����m���Tv���o�b�p��ZY���������J9o)?��8�.�V���c�PƐt
׫�J��́	P6���@���U@���:��F�6<�AT];'�2%!���Id��F.�!�KXͯ��<�ы}2�Dh��������ïI�
���͖nh���X �U:�d}�nv(�ny(�7�ͭ�s������m�D�c��QԷC��K�����@�"O�V��hoˤ���)*)�6��|P�r�����.G��~Z�7�PǨ�o*� 7�v�ԯ7�)���G�o�g��!��ZB��,�Ӏ(�˦&�-�Q^�!��ZB�;�H���o(�,ebY�sDG�\y�Ss��=�����ߗ�H���3c/��!�Iz��޹�����
���,�r�@���;c��Ǫ�'\���k͐��S ���������b�O}@���kJ�R�@�3�0so��%���[%�lM0��]{�̜�8�uW���?bS�xǠ�j�*ر��Bg��+F��%�R�X��Uq�?�f����_���¥��q!g�M6j�"Hs��a�Ҩ����r}a{���N�n[��ptpgL���_�?�d���&�M�߾ol����Rz&!Y�Xj՛���z��"��
��� �����D�2�r����/؈ъp��6?����H��efm�0z�cUL���ޤ�Y5�x�#!b�PǨ�o*� 5���Bi���eh1q�c���	?���ֽ݅u�x���|����G��8n���!#���.�h��&r��rs�(�̴Y�{'%sAX���	qn[��pt�M��.���>#���!L(��̭�d���7��a�vݝh�c�A�L'����Y�^��G��~Z�7�߼u��u��'ܑ��`Э��jz�����8]�]p�cK[��-��:�.�zΑ��$��N��E�EX�orǟD�uiM���	�f�=�er߮�r�^K������О.�����e����!�?2^�9,����_�$X�)�?����Q� Н�;@�Q�����gV��|���\j�<lG�"*���.��V)ׅ8h�{V/H��+��g&(�晅PtC�o�TI���<�jl���oJ��W�Px:'0/��v
���3ľ�Yx�<��w�怖h���X ��7��6זW��z��OQ�����gV��|���\j�<lG�"*���.��V)ׅ8PǨ�o*� 7�v�ԯ7�)���G�o�g��!��ZB��,�Ӏ(�˦&�-�Q^�!��ZB�;�H���o(�,ebY�sDG�\y�Ss��=�����ߗ�H���3c/��!�Iz��޹�����
���,�r�@���;c��Ǫ�'\���k͐��S ���������b�O}@���kJ�R�@�3�0so��%���[%�lM0��]{�̜�8�uW���?bS�xǠ�j�*ر��Bg��+F��%�R�X��Uq�?�f����_���¥��q!g�M6j�"Hs*oeu�M�V��	��y1vXD�)62�����Vc2�����Vcv�iL�D�ҕ�Q������zȐ`q�M��9�GKP�2�����Vc2�����Vc������|��3&76o��)�u����s� J������YU��Ȫǡw_��s�֙C�T&L�P ����lG�X�j�{~ ��l�j5W��	]�	�OW��F!���K�_k���+Rɨ²�a8'�(�S��D>���������!m�dM
/a�:��u~�������C�W�{vK �-o#�s�W�D)��:���
�]U Y/�੘8��?��2�ϗz�.P̐�R
{�*����_Q1d�X�f&�6s"~�T���3n���Qo�n<�!M��T�t��y��=zjm%��b�s0��R�����sF��v_}!�*("�3�\եV#�=E��r���,�Wc%�,�F�,��{��(:/�b�&�q����w~��,�F�,����1��X��WG ��m�O���Fn�\��*�J�3���y�my$�N���Uە��B�R���>_Ѩ�f?�R���dc�@z�ׅ�ؘ��N�g�c�`�9�d�L���}bg)k��Va�ir^�*�ǒړ��Q .�L��H��	W��N�g�c�`�6��X�:����R���O�_.��{Gyn��&������);�OA�uW�U��W�^�V]��}u*w�A>je`��@d3�s��(`���so6� ;h$	R*E���&�Ut�\�m�O���Fn�\��*�-�N��0:����Rl��s��R�rs�(�̴Y�{'%s�ui�铋X��q�@2F�Qx(�i��/Rl1Lk[��?�uUn���������v��L-�>Y�B��
R\��275�،��I.Ta4�>�8
j,?���z_r<E�Ԓ�WMj
D�
��Ҹ��Y�\˔t�r�W_&�����iE$A���	<M�!Euś
ʼ	ۀ7���\�����4�(r|����a�y8�n�����wNN�R�p8�<l������o�]~E1K��ꡔ @��-Y�Q-a��_��$P�_��q*�>��S��ޅ�l���3'�]�6̤뢲�
r[B1Y���zR���b���Z���21N�����D=,Ϩ4�Z\��׶��$P�_��q*-���i��1������QB�ϓzp�-a�D͢fU�9�׏�����MFi��|�3;c�<pϣ�و�9K��3̡��&Y��V�H�����-2��,���We�v����3n���4�B��ٴ���Q{s�؈9ϒ<�3z��ZΓ�Nٚ�U���ڄ�����DV,�ـ�P��>��6�����K �_��,J�l�/�D�����TeE0��WC�)�kǇ<�������y-�����Q%YD3���L����|Ӵ��^�=� �9D^�����i�Ü2>#��L_��s�֙��p���?�7r���gE�w_���g�0�u�?�I���6\�4�@���(�?<-M�O��~��D�$0�<����5>!\������dB}~�}�"R*E���&�Ut�\�m�O�����(���d��{S˥�l7%����r����1�fT_UX���-M�^���e\���6A�T��,q�����L#�>;���	ݔ�?�d���&���pP���fa��50Z��5ߧE4��p�-a�D͢fU�9�$�)�vxGY���v8N6j�"Hs:L� Q�Zm��zz<���Rk��%�.��M��	�W��ٕ����ޒ�����5�X��h�;��|B�M%>Y%�Μ=E��r����%��֊�0h�5e���a�֧�I��3��a���	)Ԭ�>@X��WG ��Ѩ�f?�R�^�*�ǒړ��Q .�L��H��	W����Ӽ�!y(t-�D��ht��g����?��ya�	�Z����(�^�G���=�ni[�b��o�CHn
V~$(|��s�i�OV��6�Ħ��spC��J��sr�l���:��KY�"橝[��+u�CX�U��w6Q,o��񐙣#�S�T�� |���t	�,^)�%�]��8��$#��pb�X��WG ��?5'[�鳥�����݄���!G����W����ref��A��y�:�B�)u�%N��x�*aE�ܸ�r��%.P̐�R
��dUb/�Hf�o7ȣ<s��X�8F�w�Q�+���z�-�z
-��|�!I/�������#�$A�X�r�J�1���K���L���4�04�jfFi��|��wØ�ߜ���,�ǰH7"LTftpϣ�و����+T"��nrm؊(����j����=���������ǝ�(�b��T�Q5<�i���(E|�����rd�d�JR'b�'=�(���?*�25����[��W�{vK �i���>oX�ȀY;2deM�|�Zi���^ =z`D�N�wv�4f��%ޓ�f�f"_qR�U�ƜzDĝ���j�3���O]�
�󑠱`�D���>��Z?�3a�.��[;T�!'tk4̑	h��[�j���-��].���=���*� ˽0?�.��L�y���4d�o|}h۰� t��]�kj�U�f��&������w�iU�c�sC�CW�[��7���̸�C�M�<4P����4�9 I�������p�<�2�Ҧ1���Z��(|��s�i�nRdd�������O,W��p��Z�SnH�B� ;��T�(�^�G��O�������(|��s�i���R������@��b#8ΓW�g��ѽ��J|�����!m�O���{Ұ�f�>��֑xGV��Ee6���uo�Mj:F�S��/�j�LY'�P�h<���8-I����c���1�ā���"�1�C��y��Π
.�a�ke[��u��}�l�1�����0���8D�K^oxkx U�_@+���Ã'�� ��,�C�����෨J	a�ЗU���HU�:=�m����y�BDG;9��Pjs��r�F([��}qn
V~$m�O���rd�d�JR'b�'=�(�q9+t�}=��Ez�wq=0�>\�(?i˸3�J�
�M�'٥��gVؠe��@F�KD�Vr[?z%CS2b�ү�+ҋ�K:+> �3�ѳ��w���<����5>�,��5�Q���1v�C�� Yz��c� ��*��؁�T^����H��	W��ү�+ҋvE7�MW��C�j�7���@��T��R��a�J��vT��N�g�c�`^��W8���'oC�XK(p��1�'\��i��ΥT�t/tyc����(t-�D��ht��g��倉r˲����ɛ�?өB�R���>_�6��X�X�ȀY;+�z�;0��`����n�Mv!���x?5'[�鳒��@��T��R��aI����Hp9��x(�i��/R8BW�R7���r_��m�d�?�4��Ǌ��i�ъ�����e���\���rK�&���&S��"��hTC�G�L奟gke�(ƚ�4j�}�������A��(/4��]G@��z"B�4��X�q�hH0��^o��[�u`���ҕ<(�(m�O����dQz^Oыq�GR�'�^�����P�HS|�4�04�jfJ�1����ݾ-/�φ��<�6�)�@����(|��s�i�nRdd�����C1zh�I�V.��S^~ߝ��wh���t��d��WԶ%T��Cz�A�uG���G�Ȧj��v������^�n��Uh�q�em�P�c`��g���;�%�L
6�,��a-;�!h^���\�}g?	��oW����
�H;"�g~����Xp/H]K�_%�0h�5e��7�b��C�����෨J	��1��X��WG ��(|��s�i�nRdd�������O�g&xdp��N�SF�e�N�|�!�������'|F��ΥT�t(|��s�i��j����F�݄����Mv!���x�e��@F�KD�Vr[?z%CS2b�ү�+ҋ�K:+> �3�ѳ��w���<����5>�,��5�Q���1v�C�� Yz��c� ��*��؁�T^����H��	W��ү�+ҋvE7�MW��C�j�7���@��T��R��a�J��vT��N�g�c�`^��W8����N�|�!�������'|Ff;[����X�H��C�j�7��s\��,��|`��=7�}|��	��a-6�Dam�O����dQz^Oыq�GR�'�^�����xȀ��D׏�����M/tyc�������so��C$WE����P$�@$�N�|�!�����a~bh?5�/tyc�����&Ř�Tٱ ���6���B�*��rd�d�JR'b�'=�(���:��KY�[b%Ɨ�m�O������W2���ݟ=�NM���ɛ�?өm�O���rd�d�JR'b�'=�(�q9+t�}Cٲ"@�l��Q�g��| �g7�ۥW׆V���m�ϣK��Z�M*x�fr���K��������I 㩓�a�8�x��^w.�����9.n�Q+��K(|��s�i���R������@��b�x�. �甑�:��KY׏�����Mrw�&�z<aSm�6��`߸��S�Ȍ3QP�B�=s�]��7�0�jv�]��-��;������l�����C�	V��΋�
,`mu��.8��l�H���{D�u�nm1�H��ۗp���x��^��W��\'�3Dm��A��s��;��Nc�4�9 I�������p���>�.?�d���&��d��L_�xw�<2%�	�}:{u�a���B�-{�=�5&��������D�$0�{���F���B
lE���Pع���a�	�+4D@=��Ez�w�W����<MN2��΢g	nܵ,�ى�1��J�b�z'hۉ)��R����\�G���Ԛ��b�$*�&�P�2�P�L��M��a�<d����C�j�7�����N��qs�p�Ehp��l[�Ƶ�-M�O��~�/tyc����s��1^~Ϩ<Z.َ�>�1O�ME�g�������(ӈ��Z��&61�\�G�����}bg)k��Va�irxֶH���k��h m�-�C��7u#md���t���(�x�H��	W��ү�+ҋ�x!!m�/ śL��ł��p|3�ޝv�@��s-�N��0�W����<MN2��΢g	nܵ,��f�K\>-h7�cL���	Ǹ�y85�{rRKC���4����U�ԝ5�c�}���F��b練J�1����ݾ-/�φ��<�6��#��.����4�磕�&�������_S1����9(�Hv|����� N��r*Ѩ�f?�R��&�������_S1����9(�Hv�($Z�u��΄x�g��	��S8�u}F�4ŕ)�y�:�B�L��X�~��LEh��� �Ne��~~@�\���0f�g'oC�XK(p��1�'\��i��ΥT�tB�R���>_?5'[��jv�]��a����g��� 75K�+���8�׏�����M�,�%�Y3�s��(`�s��1^~Ϩ<Z.َ�>�1O�M����v�Z鎬�������(����ㅣz�xHhMJ{/��1Tw��#�-�4�����8�.rɗ�-M�O��~�?5'[�鳒��@��T��R��aI����Hp9���&�������_S1����9(�Hv���D����ΥT�tB�R���>_?5'[�鳒��@��T��R��a���3,ő��Hp9���&�������_S1����9(�Hv���D��f;[���J�1����ݾ-/�φ��<�6����	��~�'oC�X(_��89�x�Վ��t�!��瀱um�O���������G%{�e���k�٩��sNV��C56j�"Hs����}=�pϣ�و����x��U�Yyr��'�al��paf��pD��x�fr���*�Ҳ��X��t-߱�~���t˛�ljv�]��'\��i�M��1Wz�t���(�x8wkd:�L'oC�XK(p��1�byQQB�v*��A9`"��T^���8wkd:�L'oC�X(_��89>�6���TZxZ@4�׻E��}"�����とu?u+��Fz���S����h}E}��3y۹+�c�	��ʤ��<+93��Cxw\8��t�1�>�z�/��-0��C���i�����K	h85>-�F`z�k��h m��.�G��:F�S��/�j�LY'N�يv����
��h�����pśL��ŴZޥ��FxZ@4�׻��Ƭd�e�Y���T�+^<�ҋ!�<�o�2JC������D�
���
?�-�Ce-X��y�:�B��=z���j
?�d���&��]��7�0�q�lN}Ot�l�1C��(�2VP��ѢKK�r��5�c�����|�\;͖�Ԍ2����:C0�C�t3Dm��A��8�iE�į��ć��Rٕ����ޒ������z��w�j�_��s�֙�����`�}�2�����_չ�ŉ�B�*����(��kkdBө��c�����|�\;͖c�M�)�v������D�S�OZ�I�u��1lz��M6� ��<;A�D��n8T �����SO�z�1�'�al��p],Aبs+��,s�3�
�=���!� �Y>�3�eZ~�B�*��Fn�\��*�T�xzG0e��w�a�k�ro��V@�Wu�t�x����T�!�J���)+�dR�L��GJOǪ;��E^���\�}g?	��oW����
�/|R-��]�����Ķ���-��ol2���a� �""y��g�0�u�i��"u��/|R-��]��A�1Wk}�aá�����-��ol2���a�H��	W��N�g�c�`��[sǱ� �Y�A?Љ'�-�����1�G��8£eՓ8���/�E�g�������(ӈ��Z��&61�ȴ��A�D�$0�#W2���j�Bd��g\�Ҳ�}�-M�O��~Ӿ9�d�L�o����Ӫ�a���B��#�fp�J�@/��r ��%�z�J���U��ǣB�Z{1@.&�<��V!���[Ѱ�^d7�v�ԯ�-�Vb� �� �Y��+�����[Ѱ�^d7�v�ԯ�`�L�i�p�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�o|k�Lb��ܐ�}ļ?E�!$6�#t�,��r��WdM4@���cꂃJ5^��7��NV�L���s =��Kݝ��+�9-�i"'���Xw�j�7���$��$@.��dR�L��G��q �2:x%�c�m1�H��ۗp���x��P�otO�OA4�*׃��҂���G� �9D^�I:�K�R)���τ��dR�L��GJOǪ;��E^���\�}g?	��oW����
�/|R-��]�����Ķ���-��ol2���a� �""y��g�0�u�i��"u��/|R-��]��A�1Wk}�aá�����-��ol2���a�H��	W��N�g�c�`��[sǱ� �Y�A?Љ'�-J�3���y�my$�N���Uە��}�u�0�_�K:+>ً�?�(�p���� L7�i��6ð��TvE7�MWO�F�Tr�f��4i�׿��/v�b~*��s�����T=7�}|��	��a-6�DaL F��j��H0;��e�B�l
��qi�տWdM4@Ȋ0�ɬ���BT�^��(�%�8�e�&���6rw�&�z<a��r����5ߧE4��p�-a�D͢fU�9�$�)�vxGY���v8N6j�"Hs�5PenWLq�"��2�BC"��`��[:���ph�9e���Rz&!Y�Xj՛���z��"��3���c�Z�~u2W��Q�k�Y���@�Wu�t��U���T:z&���qB�O[H5�Nxkx U�_@�R��9�u�1It�� ���F.�!�b!>��]H�2?k�vf;[�������,�ǰN����;�#K?�i�j%�~R�`q�=9ށ5�$Y��X�pgL���_�?�d���&�M�߾ol����Rz&!Y�Xj՛���z��"$Y��X�9<���F۪	�}a?�d���&�',+��+�lq&�3�N�0��B$���n�����9�'%��v�����X촯��c��� � �9D^�W����,��h.3I�;��|B���%���lq&�3�N�0��B$r�Ch���U=h�.�{X����O��	�����Q��m�J�
�M�٥P5���rs�i�Ǘ$� ��������,%�ۧ�A�YQ�(�O��Q�����gV��|���\j�<lG�"*���.�/��m:~Ns����8�����������'���Xw�j�7��5�K���(~N�[��F�r�f�t!L(��̭�d���7��a�vݝh�c�A�L'����Y�^��G��~Z�7�߼u��u��'ܑ��`Э��jz�����8]�]p�cK[��-��:�.�zΑ��$��N��E�EX�orǟD�uiM���	�f�=�er߮�r�^K������О.�����e����!�?2^�9,����_�$X�)�?����Q� Н�;@�Q�����gV��|���\j�<lG�"*���.�/��m:h�{V/H��+��g&(�晅PtC�o�TI���<�jl���oJ��W�Px:'0/��v
���3ľ�Yx�<��w�怖h���X ��7��6זW��z��OQ�����gV��|���\j�<lG�"*���.�/��m:PǨ�o*� 7�v�ԯ7�)���G�o�g��!��ZB��,�Ӏ(�˦&�-�Q^�!��ZB�;�H���o(�,ebY�sDG�\y�Ss��=�����ߗ�H���3c/��!�Iz��޹�����
���,�r�@���;c��Ǫ�'\���k͐��S ���������b�O}@���kJ�R�@�3�0so��%���[%�lM0��]{�̜�8�uW���?bS�xǠ�j�*ر��Bg��+F��%�R�X��Uq�?�f����_���¥���锴�;��|B4Y-<L'��s��;��NcQx�Ԏi���QQ�W��vw<&?������Z���Q��m�Ү����,j�W�q�l0���2�W�ub���<p�ve�}��i�Ɣi�����Q�@�p�~ge?�΄x�g��	��S8�8�{�G�ÂJ"�Kv*���V)ׅ8߼u��u��'ܑ��`Э��������'���Xw�j�7��5�K���(~N�[��F�r�f�t!L(��̭�d���7��a�vݝh�c�A�L'����Y�^��G��~Z�7�߼u��u��'ܑ��`Э��jz�����8]�]p�cK[��-��:�.�zΑ��$��N��E�EX�orǟD�uiM���	�f�=�er߮�r�^K������О.�����e����!�?2^�9,����_�$X�)�?����Q� Н�;@�Q�����gV��|���\j�<lG�"*���.�/��m:KXͯ��<�, �dh��X+)%`d�Y��ïI�
���͖nh���X �U:�d}�nv(�ny(�7�ͭ�s������m�D�c��QԷC��K�����@�"O�V��hoˤ���)*)�6��|P�r�����.G��~Z�7�KXͯ��<<qJ�A	D�0��E|�,�Y���҇�d��Lԗ�'r����MM
��,=�����yU[I���W���'h̟K.�0�N?c�<��6��ߗ�H���3c/��!�eY�r� ��[O�"��!��ZB�;�H���o�#m[)����6L<aMYߍ�?`غ��φc��5p����U�:�	��0i�wן�
��0��᭖K��"h��3c/��!���z{J�۞h�G��D9�{w��Q��D�w�����h4c�Ү@;���! n@�����!��ZB�d��Ꞌ�kL>�`��Ee�&��c����[�����@[�_zβr�v��������Q>�^2�����Vc2�����Vc2�����Vcl��w&� ��tF��J�����{��ܨ���[����9�GKP�2�����Vc2�����Vc2�����VcSd�*-}Q��eh��2B�k�`�?��<��j�3����ǟ�u�o�e�d�`�n3ԛ̿b��Y�PG�(C�A<�Z��B�\��G�8�*�# ������a�<^�>�rK�r���a��HlQ/��?HY�S�h���f�w��)�@���*�nӜ��Hǈ)T�u9���3;5��ؙjl.��{
��m	���Ʉ��:�5[�] �4�$F��߽��tQ46- 	Iz~�Gy�'W��	]�	r"Dd���꺖Z(��!�Q���y�,n���w�� ��5�AkTRY]���p��1�����+?��5b��Vu���|/���ϣ[���A�*w!�I��=� I	y5z��<$�W��xl��2g���z`Ε�ھ�i�䰥�R<���Jq���x�t������5���֡�&Y��V��O"�|:�@���*�n���W����]�lEGV`2ɬc��WN<�V�QK�}2r��q
�T�P�y�'�X�6q���D��$B�����o�u�/|�Rc��[�jZ���R\h�(E�4��+5��N��M��q\�!P���b6:Z��c/����1m[�d��%^� r��DI6�<�k�`�?��<�G��-^/�eo�L���hl��h&�.���Fٷ�p"�.��탯;\߰{�P�1|j�:"��8ļ���N}�O̡��Xd!����y�8Tc�A�Gd�o[b*7+���Ã  i�aT�V!��;fcMy�KX��ikj����ے=7�}|��	D��X�*��_?�v��9�2�L%J�bb��|;�����8������t���MIV��8Y��I/��\]�3�� �frw�ܲ��}([��}qn
V~$���ȏ��F�[�c�Ĭ	�g����#k�˟ܒ�o|k�Lb�5ߧE4��J�1���k_���b_!2�͞nOY{�q�O� 	�m)~�l�wv���f��U;ߟ�+�X`��_/z��w���*#�IQ܋��5&��J�(�딻����/|R-��]�����Ķ�(�^�G��%���}Mv���-x��p�̼�d��Ꞌ6?
-9aƬ��;�Ӏ׬�����D�{�I`�	-�_3�mE�_s�rp� �1x�it���w~��,�F�,����1��X��WG ���zt��[��t9��\�w�xo�A�\�G���o����Ӫȸt���(�x�H��	W��.3��؁���Si��i�Pع���a�	�+4D@��~JFNǭ_����頴��j�n�q�[��9�Χ�˓#����<T���&�jW� ���_(�a�x(�i��/R�������	սL��$��R��	π2�����Vc2�����Vc2�����Vc�1�^A��+��,s�3C[k:!L)�e�C�$2�����Vc2�����Vc2�����Vc͞���� pbL���(�q6?��O�z�`Ɵo��FZ��ժ��*#�IQ܋
�:\߮��+r�mt_��'��A4�O>J`��dZ0o�vʺ?�ο�\�#_L��
�xw�<2%�3o� �� N��r*M`B�Ӑ�W ���t�-M�O��~���9 �v�n�������%��v�ښ �{��{Ѩ�f?�R����_��
�Q�Xn�)��d��X��WG ���i��"u��/|R-��]��A�1Wk@/��r �a�<d���T�����݄���'٥��gVؠe��@l�ްX@�l"�p��^�F=E+=7�}|��	��a-6�Da��q�GH#����N=f;[���J�1����ݾ-/�uu��ڿ׏�����M��ܐ�}ċ�PkO�׸`49�<g?�U~a��O��`�`Ƅ.�R�+9Gì��W�'�,|�M*����97�v�ԯ硙�t�\#t�,��r��WdM4@�4gՇ�*�� $)�lj�iE�EYZ/�VU�簦-�b�+�