��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-?H)t� �hz2��ƿ� �lJE�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hp���Ť�Mn��X)r����#�L������5N�1 T�V	�tL��	F����1��]}|��~����S˶���
>�1FaO�.Jd#$f���|����yRu$k��R�9�#��f�mX����$[��`M��
�k �p&II���<7����SeN�7��n_Kǈ�V�MT7xB2I�d�ߟ��+�+�n��po�>g1�]l�&Y��F}갨y����K	����2z2��ƿ� �lJE�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�iJ[�FUԥ%���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�ħƿ�9c�1��8�h����,����^�V�.u'a�zHF�$���خ�q>?�=�T�x�JYI��'��.��y7�N�	O����[�i~��'n�^0oZt�Op�t��5����`K�wN�3�d�����}zES���)U{݇��*�'n�^0o�m�0Q�M��5����`K�wN�3�d�����}�11��Sca�&'�'n�^0o _xB�I��'��.��y7�N��b��%��4e�w��~tR6�\�zL͊�q����#���1�o�$C�,ݷ�:���B�c�`a��T��w~tR6�\�zL͊�q��QX~�mrHO��c�Y01�������Vz^�Y�uzL͊�q���t��m��RK�F��ޯ��E����T��IC܈�,y�,�����D�1���LI�.�FU���A�"Z鎬�������(����fS�X��C�GI$��ǂcY�~遅��'�:��'n�^0o��S��S�Ib���ό���.ӭ��L���r�Ͷ�7	��4�kC2�_����*_pר&Vv�'n�^0ow�?�b�>޼�\�v�GM
�-��q�N�ܔ�L+�b�?.݁ei���J\��g9$^>��U�:/��<�W�C%���80�va�{����_�=WB�'
Ү��p7��e�1Eu�J���"�8<�V�Zs�f�f_G�_�(,/;���(�!�q����e+X���.�b�E�<�W�C%q���B��<�W�C%���80�va�{����2��� ��b�FP&
�c�,�%Ah�%4
>��XP���/e��IƬ!��Tӧ~�k�X��WG �����n�O�V[���yuj}��8�,�[�1��}�x(�i��/R�9��o�����Pm�TT7���1���|�@TߟW�����m�ʃh�[�x�o�~�<�~�V6$়@�|�\��9$����:������ț{@�P}��O��^��mi9�g#���k8�<4 ���3�ҺIÙ=�H
,�L�F��KX��ik8X:Dn2(�-M�O��~��Z>H@��L��>��B�R���>_�Z>H@���X~�� �4�04�jf�y�"�V���Ά��߼
�d#�sBQі�㖏��ś��޾&�-��)���p������8<�V�Zs�f�f_G�_l���P�/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'���?���ʢS����E@�ޗ9(����	�^��i�ħƿ�9c�J9�^c�5������Փ��ખR���=ە���oH��O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���[�}c��G+�
�c�~R;}��I��1 T�V	�tL��	f�g���Z�ʣ���xMf�TS=&��>�2���pM�i��w`�1�B�G"��������K���!z����vYvI�͌.�hMR�`6�6p�����w�vln��������7���*�����;�(i^�0�|�U�L�2 �Q[TH���"�,�>E����P�1�,�3�T;���n�s��?B�OWF��j��
��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����@Kprd�t@0�
y^ �\#+��S�M͈�{�P��j.Z��$�sӢ�]3�����c��(rKg!�h��� $��:c+�I���y���OJHn��z���G7���� $����oa��ܛ�	���������IÙ=�H\[�*H'nLѠzM8%�Y~��`�JKݗZ:���'n�^0o����y�]�\�۟�-?�d���&����{ԕ�h7�{`��������K~�5N��
_�,|��7�On�AN�.7����,�R�A��%��Nt�ꬡ��k�*ί��Oi��!�`�(i3x�]�V����:L��:���H�����_n���!�`�(i3!�`�(i3l0��F��j �i7�sp>��cg�ų��'�oD�!�`�(i3�Q�^�y�zL͊�q��[�į��OƋ.]$�����m�!�`�(i3JHn��z��r9�3���Z8"�|o	���=l!�`�(i3��Q]� _�rs�i���l?��	D�ǲ�a��x����̄y�����!�`�(i3�n`5�fK��0z�cUL�ӒN��G�/"��]�Ͻ!���<��!���<��!���<�AF9��ԸS~V]Ŧ�^&�c��J""�,�>E����\�vūx`��:�͗}��Eނׁ�4^~#h=y��l0��F��jT�����N��'�-qNↂ`Z"�Au,���Ex��#��LzL͊�q����UI�hI<a�F0�-�?@���w 񕮘K{BJHn��z��r9�3��y��p>�R�/�]Y`�!�`�(i3���+�J��Y�{'%s��.|Z����=�Q����-���+^�V]��}��ł�!r�dN�<@Iv��nt=:���S��Aj�X����~Y�({���K%J�"�5M�U�=��<酀�ʭ����@�)zL͊�q���[��:�
*�&&_E�P��$�V�)���N�N�F�39���XP���V|����@�Nt�	��um�L��$k���[	щA�b9���:&�>��s̬���	p\���z�4e�[U���z{�w�?[8T���`�v���Ŧl<�8 v�>���|!t�נ&�_!�`�(i3�E����F�'n�^0o����y�]�{�6�e�]h�����!�`�(i3�b9���:&�>��s�{�b1乌k���x�]�V����4�ʛ9�����	�����o3�|05���b����qhrp@�����7��V\s��z ⑉^_�����S#{���>���9��+�����I�Gn�V��vKn3g�)��C�+��1����Ƒ�$N�������쭯�J$�;P��� 5eI�9��&Y|�M�
!ǥk�}�`:��Q1!�`�(i3JHn��z�|=8�E<��FzBR)��p���̈́EX���MD6:�z��e,���� I�N���������)<��CB-]�;���c�`�q~�l)�������5	��]�!��vH�/ӟjZ����R]N�By3��<Z鎬�����;L�=Q�<1(f}ظ6��d#(-�+xk^���1!u7}:N�By3��<Z鎬���������k�^�d��d}7Ê7�E�4'���Xw/���:;aR[�T�.�W���1�.��eȱ�9�t�5ńҋX����|P�������A�=�8bH���L��B��K�-)K�7Ê7�E�4'���Xw/���:;aR[�T�.�W���1�<�_9���� ��H�Q�ҋX����|P�������A�=�8bH���L��B��o�fy7Ê7�E�4'���Xw/���:;aR[�T�.�W���1��~�yD݃e>���K�l�5��E-&�1d�������E��@IE�U��@�ڗe'9�C�،���S������-��uO����(�{��{�{l�f|��rs�i��)��7���n�EdF$�c|��)�ȣ�uB[U ��̇�ji�yHe�枘#�a(􆿳�i�n����L+�b�?.݁ei���J\��g9$^@"P�
BO{[���G��D�P�E6�)u�ҵ��B@����������5	��]�!��	Ǹ�y85����[��3&��㖏��ś��޾&�\����W�G81���5�oC?�Q䨈y߉�m�$���=/�Y%T��BPS�)37J*uc�A�L'�T��ݙC�a�	�!��g��U��\�e��)��E�>4p���eq��$�'	��hyﭡ�����A�b�*܋���ԓ�Dd�3�[i�`#�Vao�r�̏[��v�$�(Ktk��^h=g�^)�I��w��,����Ȥ�(Ktk��^���ֶ�I��w��,����Ȥ����I8�h�"B��$I��w��,����Ȥ�JT_��
�����I��w��,c�A�L'P���6��G�C��Y�K�za۬���f��yd�x�RFgI� �8���:�k�ay�k
��{�#sc|��)�ȣ�uB[U ��̇�ji�yHOƋ.]$�6�7��8���/�A���0v7���V�x�O`�����
L'���Xw�j�7���$�� %X�|����OC��:�|.���u*�c���E�?G��g��U-�e�M-n����w�o�FAMsYl���#�]�!��N��7|5�dH�M�$/Yl���#�]�!��N��7|5�Y0R�ne�Yl���#�]�!��k��v�Kp��}�G�@����uO����(�J2)V��(�
t�ژq���U�$��	�fѥ�[���В����m8�{w�d �������E��@IE�U��|P�������A�=�8bH���sA���U%���;$��]2�y�Z鎬����L�`u�K�˱�Ui��Q�xy}���
Ч�P�2ݙ�TD��-�`��8�4�%��mz%���=a\�&'UR�q���t��	�dS\Z�vm������SJ��8�CW��Y^�i���,�qm�c�,�[`�/S�B���7G#+��Q2�+�Yɶ��,�qm�c�,�[`�R�l6j�s-7G#+��Q2�+�Yɶ��,�qm�c�,�[`���T��S=�7G#+��Q2�+�Yɶ��,�qm�c�,�[`��Ak��_7G#+��Q2�+�Yɶ��,�qm�c�,�[`�Id����x�7G#+��Q2�+�Yɶ��,�qm�c�,�[`�A;s���y7G#+��Q2�+�Yɶ��,�qm�c�,�[`�-r__A)C7G#+��Q2�+�Yɶ��,�qm�c�,�[`��Zqx�٣7G#+��Q2�+�Yɶ��,�qm�c�,�[`�������n�7G#+��Q2�+�Yɶ��,�qm�c�,�[`�Q���47G#+��Q2�+�Yɶ��,�qm�c�,�[`��p�����7G#+��Q2�+�Yɶ��,�qm�c�,�[`��x�הsD�7G#+��Q2�+�Yɶ��,�qm�c�,�[`�c�-Ϗ7G#+��Q2�+�Yɶ��,�qm�c�,�[`�I{�i-m(�7G#+��Q2�+�Yɶ��,�qm�c�,�[`�H�����77G#+��Q2�+�Yɶ��,�qm�c�,�[`�e=��Lx-;7G#+��Q2�+�Y��Fi4NE��<^&!!HYk��\�*]ݿi��H�4?"���і�t���,���5��Ȣ�{l�f|��rs�i��)��7���n�EdF$�c|��)�ȣ�uB[U ��y�~ J�~��3�@[��
<ݓ�y���õ��Mn�k
��{�#sc|��)�ȣ�uB[U ���rШ1�ץ"�m���rD�P�E6�-�4,�#���7|�
��(�
t��Y�{'%s9j�G ����.Y��㖏��ś��޾&�\����W�G��#*<\}y*�����T�\ ��q��<P�Ϯ��㖏��ś��޾&�\����W�G�{�6�e���=���
�'i�! ]���f��v�鳔�Ċ��8���K(��z�j�;9�e��L53����+��V�W�S�w҄�+�va��2��Ft
X�&��$�B�I:׷�Fi�k�Zׇ	JHn��z��k"����_<mDrW�B��ɥ����%�a�HL����rm��U}�	w�v�����zL͊�q���zH���u���oa��ܛ�	���8z���,�v���.�/'��Y�
JHn��z��k"����_i��Rp�������О.abK��W�󕏜9����Ÿb�6���.c9_��X����w$���ｻ�b9����^����$���ｻ��C��J�cu�q��]N���r���L�\��N�[�}��|�}�/U��`A����X�Z���#I��'���k�8�]!?늘�?P�v�
���"�m���r�b9������kR\�~���ێ`*Q�UK�A��Ujy�/5;�Rw���.h���S��9�[vĄ4Ȝ"nF^����˽�ْl��]�B�M:��2�R�)��<|�9�a��!�`�(i37�ܥ��2������\#O���o��z>�n�SSC�	��X�6X���(��O��ɀ"���Q�^�y�����9�!�`�(i3�yw���-��C�	�v��Ŧ�2ެ�x_/�Z�s��C\����nh �C�x�Qkgw��.�޹B$~s%��@�:���7s�o~U��A��C!�`�(i3�Q�^�y����W5k���(�8�t���wM/�;z5�z�Hf�!�`�(i3 ���3�Һ����R-�,JQ���q7#�nbk*�,��!�`�(i3%Ah�%4
>������GޖW�/�
�^�=�Q��M:��2�P`��dpfV�L��nw�4��P�vzo��f�(��q��P�� ��S
e���z��P��J2)V�o��C!T*�q���U��}_v�P�ڜ;�
_���F�-XX!iY%T��BPS�)37J*u)T{6T'� ��S
e�CHD�u6�ys�yze�Zv�o��C!T*�q���U��}_v�P�ڜ;�
_��q�X�Y%T��BPS�)37J*u��xc�l��m
��5�(����r��9]�Y(R�_�'O��~E=�I�t�5ńҋX����|P�������A�=�8bH����@�]���N�� Ќ�}��()���V�(^��<��z��}�����z����A�b�*܋����؝w��p8� �`e~�Ԡ�i�]'<���RP=	P��{l�f|�-�`��8�4�%��mz%���=a\��J���� ��S
e�CHD�u6�y�=���j�9�o��C!T*�q���U�$��	�fѥ�[���В����m8�{�X��R��oC�z�C��^�j��Ř]2�y�Z鎬����	�+9��\dn�'c�����ze�@�!����8�j�.F����=	���3!�`�(i3��{l�f|��rs�i���1L��I�G�C��Y�K�za۬���f��yd�x�9�K�^0r߼u��u���T�\ �͝�����uw&jt����&`�?ӄ'yy*�be�C�8�%��"B��$I��w��,c�A�L'�T��ݙC�a�	�!��g��U��\�e��)��E�>4-���*(߼u��u���T�\ �͘�f��p�b�z'hۉ)�$q&PbOG�p0>���h���R�a�R����G=X��P`��dpfVW���x�Ai�_,+2����J.h�&�0`yS2|�Z�F_u�E����F7G#+��Q2�+�Yɵ�Q�}�qjZ����R]Yl���#�]�!��U(<�i�uwd�ч@�.;�<.��(�
t�ژq���U�m?��q�X������E��@IE�U��|P�������A�=�8bH���cN�Z�3J��4��>j�5�i ��TD��-�`��8�4�%��mz%���=a\��J���d����(N�̴K��U֬����
L'���Xw/���:;aR[�T�.�W���1��gt�k�T�^��	�Yl���#�]�!��k��v�Kp��}�G�@���m?��]�b��ގ�2�	Q�o@IE�U��|P�������A�=�8bH���cN�Z�3��b�ђ�3稨�;�<��z��}�
��|�6|�+�� VU+I��X��8����]K�I[K'�/�ޑf�������~T���١��yퟻ�xʸ�fْl��]�BWa9t���V�\�۟�-?�d���&����{ԕ�h7�{`���@�	��h;E����<mDrW�B�����W�^ֻ����XP���"Ru2:#<mDrW�B���BC?T�vx�#ã���\�v�:����`Ё���=�ɤ�c�PƐt
׫�J��q{�f��a�:&�>��sAj %�Ho�-[�v:v�o���+����7X��U�?	r��;C�(�oR�)��<|�9�a��!�`�(i37�ܥ��2�CH�(���r;��*!�`�(i3"�,�>E����\�vŘ�xQG��tp�p}!�`�(i3�E����F�_�����e��[]qE�&���W����Q�^�y�N��B�)YZ��ͨ�(ͻ[$��6!�`�(i3���+�J��Y�{'%s��;d�����M!1�"�el[��� 񕮘K{B ���3�Һ�j_ R�ϴᏅN~z��9�{�G�K*V׹ږ��_�(_�<���y���2�&���	/]�����F�>l0��F��j�4"�I<a�.��y7�N��:�h�!�`�(i37s�9���o��S8��#�1e���d�Z�O����	a(􆿳�tP"7��%e��0�U+�qbp@�
\�`�x]��n���B>X��
 ���3�Һ�j_ R��<�Pfh��$�o�]��y�߀�����Z���<�a������!��٫����y�8�>W��M:��2���,��]�x�ze����^Eѫ�@���;)�nrm؊(��v�N��!��c�e"_�{�qЧǒ�E����F�ҋX����@�ڗe'�@
l%��E����F�ҋX����@�ڗe'�U�� ���r��DB�����Iq	��u�.;�<.��{l�f|�ό���.�q	��u���(�a�肢�{l�f|�-�`��8�4�%��mz%���=a\��J���5��ܴ>�Y%T��BPS�)37J*u��xc�l��m
��5�(����K�ZZ���[�K�-)K�7Ê7�E�4'���Xw/���:;aR[�T�.�W���1��8�����{r �<��z��}�����z����A�b�*܋����)�g����I(ީ��Ųo  ��]�!��k��v�Kp��}�G�@����9��4�ьb2up,�Ҹ��$��S���O��\r���㯄�����
L'���Xw�C��!a�<1(f}ظ6��d#(-o秾�!(�K�����b@T��ҋX������S8��� ��Lu�=wxk�ay���K�)�P��|�b�@a(􆿳�e�&���6@�[,E`tY%T��BPS�)37J*uc�A�L'�1�d��.�e+X�&3y߉�m�$(�K����Ο]_�ҋX������S8��<��Qʵ�'t��t�W��hyﭡ�����A�b�*܋���ԓ�Dd�����3���R����o秾�!c,?%�J��l�� �7G#+��Q2�+�Y�RiP���uV"��J���TD��ό���.�tl��(Urs�yze�Zv��(�
t�ژq���U��;�j[������V�p�����
L'���XwqX̀Wڪu�a��	e�.�e+X�&3��%�%��$]�6���p��HM�e��`y����;�j[�����V�x�O`�����
L'���Xw�j�7���rcJ]�0ݫ���Uh1�+\�41��w�o�FAMsYl���#�]�!����[��0���a�D�"B��$I��w��,)T{6T'�3�Y�� g�C0�C@IE�U��|P�������A�=�8bH�����m�m�&�}!$ �Yl���#�]�!��k��v�Kp��}�G�@����;�j[����K�-)Kڬ����
L'���Xw/���:;aR[�T�.�W���1��;2Ϳ��u;�RH���TD��-�`��8�4�%��mz%���=a\��J������15�-x�B�G@IE�U��|P�������A�=�8bH��Ę媌�+<�,E9|.���%�S��v���?�R����o秾�!���,�qm�c�,�[`�/S�B���7G#+��Q2�+�Y��J���۞h�G�R�����u�TD��ό���.�tl��(Ur�f�;�>)��-��Zz����(�
t�ژq���U��;�j[���K��e�Igg�QuU���������
L'���Xw��U4�i�PG{��_�`��B�0w��]2�y�Z鎬�����Vk$Gɶ��'�SS���L-�yC³��O��!�]�!����[�����2��C}Lr<[�M���h�$I��w��,)T{6T'rF)���X�3c/��!��8�ۦ@IE�U��@�ڗe'���,�qm�c�,�[`�������n�7G#+��Q2�+�Y��J���۞h�G�rv�Bj���TD��ό���.�tl��(Ur�f�;�>)�Ĉ��^A��(�
t�ژq���U��;�j[���K��e�Igg�Iy��A������
L'���Xw��U4�i�PG{��_����c|�	.Y9��O؎QZ鎬�����Vk$Gɶ��'�SS��/ل�� �CX��V[��]�!����[�����2�����ǈݻՑ���"�sI��w��,)T{6T'rF)���X�3c/��!���L���@IE�U��@�ڗe'�;�x������d�kⲘ�]��9^�)�l��j��~+�����dh��TD���rs�i�jw��k�DUK�A��Ujy�/5;���"X��[�`�L�i�
j��qZ1D���>.%d�ҋX������S8�@~m)�/�e���{��T���:F�X?�g��U-�e�8JH��ig7���c��;e�0
A�����)��䀌�yHJJ�5H��z���8�ǮD��ߡ(5��d9`�v�����襰(���qN\r��`U(�M�z���N�?��]�b�r��o��C!T*Y�{'%s���䒼���Ÿb�6���.c9_��X����w$���ｻս���`U`�4m�T�4��r:��
����m�G\O�E朦�T�\ �͍��,dE��'�ƒ�s v�H?��B�٘�N�?�����3�ht�����
L'���Xw�j�7����k�8�]!?늘�~M�p��=�hXV��C$��	��c�iUW��AR��C�t3���lR�1屖ʨg��U-�e������!HNi�֌� �����mƮ�ʰZ�	��D܂�A��W8ƭ��K�Q0fߛn�xSbI���Z鎬�������(�����ݬ�g#�)���8����S(�{�6�e�O
�_�Z)Z�n��[��{_8�Y��=�}�Vݨa'�<� \�H�f��X.sB��ÚT����/�!�rs�i��UQA$�|x�5c�@���v�8:��$���:F�X?�g��U-�ee�@Rv����my$�N�����X8���K�Q����D<&�V����S�d�٣��c�A�L'k.4�7�Ok�iUW��AR��C�r`$ܧ�T�����|x�5c�@���v�8:��$�ıxJ�P�a(􆿳�tP"7��%e��0�U+�qbp@���K�Qhz`��I>����}ge�d�٣��c�A�L'k.4�7�Ok�iUW��AR��C�r`$ܧ�T�����|x�5c�@���v�8:��$�ıxJ�P�a(􆿳�tP"7��%e��0�U+�qbp@�pzl��a�N����|�`�٨�U
��XC�d�hq'���Xw�j�7���$�� %X�|����OC��:�|.��xh��M�t���&�g��U-�ee�@Rv����my$�N���Uە��ݓ��E������F�R�I��A�����J�\�)��'���Xw�j�7���$�� %X�|����OC��:�|.��xh��M�t���&�g��U-�ee�@Rv����my$�N���Uە��pzl��a�2)�,���Y^�d��d}�n`5�fK�Q2�+�Yɳ
�CӞD3~L�uIş��Y�����d�٣�����6>��h�k/���;���ͳI�E����FZ鎬����Y�V��#q>����/�����	�����+�J���q���U�$��	�fѥ�[���ВZD���zQ8���L�J��4��>j�5�i ��]�!��k��v�Kp��}�G�@���pzl��a�\���	��6�K�-)K��n`5�fK�����z����A�b�*܋���QOr��	}(9G�t/�o=�<*��Z.��0�W'���Xw/���:;aR[�T�.�W���1��
�CӞDat��ʲ��+�L�)�{�d�٣����xc�l��m
��5�(����3�Jp�����[������0It���Q]� _ό���.�QK�>;?��Ϥk�;��|B}ø��y�w���H1��@�	��h`����Y-��J��׍���ebCb��Q�-�=p���BC?T�׷eh��S�֋��8�	x�9�E�\����8�i�`!31u-��`��E��ɧ���7�)a���%}D������h�br���lpda���\��6m��B��${��?�J�Z��]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gV��Vv;�Oe�d�#���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���))~�� ��-[�v:v�o���+����7X��U�?	r������fD�!l��Q�POR�~�icҦw�xۡB;�����+,r*D'�|8܉-`�6�zZ��۸9x�z���i�>R-Zx�ItL�5�5z��eU��m�H4�c���-/��S������[C������l��WV�#a�_�ŃJ?k�mv��}0�-��D!����ހ��g�R��%ȣ��.���E/S_��c��^�
E�3���7���i��fj9�[vĄ4Ȝ"nF^����˽�orǟD�uiM���	�fvM щk�̬���k�*ί��Oi��!�`�(i3/�R�3�ݏ��A�D�īZsٸS~V]Ŧ�^&�c��J"�&8�,�6�[S�?��)(�"�}$�1=���iGn�بpp		���@!�`�(i3X�PC!$�؁��wM/�;z5�z�Hf�!�`�(i3����+��c�"�m���r��I2�	��1�7F0��2�&8�,�gЯ4H]J�bk*�,����l��;�4~���;A����z��Bo���+�ހ��g�R�]��-5L�-0���+�A6#�a)*t8l��k���ڜ;�
_��j�;\E����X;p`�#�$���C[ g��L(R�_�'��6��I�g-��&1f9m�҃��OO�!�N�� Ќ�z���O���[���U?}Da��%t�f��k�'� �`e~�����.Ԭ�(�a��c�X��1[�C�ߌ� ��S
e�CHD�u6�y�
���t�n'�Wzp1�4�����:ܲk3�� ?9<��WI5�տ�G�9w{��P�o����T���\�H_�����H���JLc�Ո�D2�^�7��߅Lc�Ո�D2��OO�!�N�� Ќ�5M�N�]�od���Aь��8#���#�����q�k3�� ?9<��WI5��0It�w{��P�o�+b���#�,�%�Y*m�/��!�`�(i3!�`�(i3:����q�G�k�kW�P�\BU@�PWMv�G�nDy��kƱ�
M!�`�(i3�X;p`���AZ�yBwV���x��\�C���K	PZ�
6�,�%�YP`��dpfVW���x�Ai�_,+2����J.h���B*y_�ϱ��[��f�8T��<�O�m ̾ie?���2|��xE�%ıν�D���K^�)3~L�uIŮ��Wӭ�6d����(Ns�yze�ZvP]c�a��ʆ|�3��8$�*�J��s0P_!-��\���	��6�> ������gt�k�T�8?�H��������ceJ��4���A�0sFw�d����(N�̴K��U�P]c�a���U�< `-�8$�*�J���A�.�p=qW�e6!\���	��6���^rg��s ���/i�]�b��ގ`ڱR̒d����(N��@Wk-ɢs ���/i�&�1d���X;p`�d����(N��r��6i��RN�-#�����E�F%[j���y㑤3���S>���[!��4�~$���'��֥���m�/��h�P�������i��fj9�[vĄ4șvU�ɹ�L�,\ަ�It}�0�.�,}���wQp��O��S�7�A\(�+�D����k�*��	���԰�I#��t˧D	��t�a�Q�DW�좘��o�$����jݵS'��㎹�a���ѳ2�?���C0�*�Y��'�oD�N Wڰ��
/Üy�a
�����7��F x>H�|����SU����o_������)�ye+��W�Oae���/"�O߸�S$��£��v��m@'�V��E�;��k�7V�<1�Mb��\�γE�;��k�7����b�Ѱ>r;𜐆�`Z"�Au,���ExpL8������l	m�� ���G�����k��k|�5�9�<�ɪ0<a�F0�-�?@���w,�6��c9���M���gB?����3�����4���`6���k�{*K�X�*�܁鹨�`6�
J1!��]c�?1�4�N�#���E6�h�+]kQ|� ��gЯ4H]J�bk*�,����l��;�4~���;A����z��x�y�k��(�a����<��j(��������J��Sծ��[�$P]c�a�����"�_�G=X�����W��y�-��\���	��6�pb|�@�Џ�F��f�8T��k�b��!�.�|Ћz�*���r���ȍ�)0f��
!I���k�Ӟ5��������Z��K�-)K�_�I�6�k_N j�S�,ċ͸�O?�^��	������ce��JԶ�.�I��$��)$磨'����τ�\���	��6`���P������Z�^�j���_�I�6�k_�����TDW�S/f��e	'�����wL	[]��$'i��7�w7Wp-��(����/��*��8�,wO��~��mL�+1���K��N��9p-��(����/��*	'��K뀚�1�]��$'i���/��;p-��(����/��*RiP���uV�Q(��r�{	u0�zL�~�'Vb�l����d�v�c�����p�8�٬v�c������ � ��<�K�k��BBI��?0�q�(� l����d���V�p��p�8�٧i�LG0�g�o�3��ҝ�b���l����d��V�x�O`��p�8��&1f����g�o�3��ҝ�b���l����dx��������p�8�ٽ0�.&7�M��
��|hU�c���姻������vP����I=[.4���^we�I��=���A�0sFw�G��mO.��X;p`�G��mO.���� � ���G�8�BBI��?0�*o�W5rl����d�)�ޭ-���p�8�ٍ��^rg��l����d�o�fy��p�8��`���P��G=X��<�,E9|.���%�S��v���?�R����o秾�!�J���۞h�G���HY�� ���<��S�۞h�G��"j�ՏDtl��(Ur�f�;�>)���{��Z�����]h�f�;�>)�|[�t�3�l����dK��e�Igg d���U�d��p�8��K��e�Igg d���U�d��� � �'�SS��[%�lM0���儘^���'�SS��[%�lM0�D"-�(�>���2��h"r���3߇�q_���2��h"r��f��k�-rF)���X�3c/��!+�d��rF)���X�3c/��!����L����J���۞h�G�]8e��Q���<��S�۞h�G�$U��'v��tl��(Ur�f�;�>)�k`�+Y�r������]h�f�;�>)�C~2�)0I�>�ܖ�4��PG{��_��9z�AR�w�>�Z�'�PG{��_��9z�AR���� � �'�SS��I?�KǶT��=k/#��'�SS��I?�KǶT����#�e�rF)���X�3c/��!7bIEH��SrF)���X�3c/��!���g��綧�,�qm�c�,�[`���<{fʹ�k�m���c�,�[`�eZ�ۿ1��J���۞h�G��${Om<����<��S�۞h�G��5G���mZl����dK��e�IggI]eLu���p�8��K��e�Igg�m����>�ܖ�4��PG{��_����S�]p�~�W�û�PG{��_����S�]D"-�(�>���2����I�}jL��s�w�����2����I�}j�I�޶Sx��2�D4 >V�`b<�.�$4����B�P�{صUK�A��Ujy�/5;���"X��[֗Q"t���'Y���,=x�q㞒��\ɬg��sB��ÚT�r��*!K�>�Ō(_Ma�~�Ǔ8���/���(M���9��m����e?�d���&�>��3�x�2I�Fq�Y�vL���5�����~��"��q��t�Pr�d[S�/W����xm�O� 6�/Y��|8�����ˏ����J*��Q��B:���o��f?~�Q��\@
����4j�;��|B���	�I��/t���SXe�Huṟ�5eI�9��&k+8_Џ��"�֙"W�}v�wO������oX �5�D�;E���y+�-���vl^:�"�P��SM*)��g>ɟ�h���B� ��~��	�c�4�b���	}�@�x��JI� ºdR={H�3)-�vL��|�`�٨�U
���9D����Q��m�4mL���n���"�A�Y1$0ZG��n�C���T!v�G�nDy��9�k��ߑ�`��å�X@��/k��A"L<hfb�{�>�v������F�R�I��A�����L3�)�oŻ�&ǥ�̻����.���ܐ�}�S��/:+�e6j�"Hs`ÀB L~��^V������_�&3� �iY��yQ=Ԗ/­�`N�(��Qx�Ԏi�$���ｻ
�HYF�@��H*����&���	/]6]����e��Q`P��^���\�}fX�
�61��*ތJe�*�O&�Wd�L�O�i�N1��!�;������^k)ٶ�m�R~�k_3�o_����M�!بDL�[��!y��Ȑ�4�(@�Q���Z��a���M6��f���}�T1�XK2/��������"�,1N��2�t�9)�.�$4���s�IH}�F[�t
�d��EZ���ފ!|�$��K�����.�$4��Ŗ��3�ht
��W�$:�-�Vb� ��.��y7�Nh�V�4��G C��0k�2�gŜn��VS:�khךSi/[��"��?u�F��%��>�g��U-�e��?���s��ʟ0B>���{��xA!P�~uQ��)�m��
e$5�
m����TԒ�@r�ADs�lE��8���/���R���7����X�l�eo�s:�r�,�n�c*$�7��c�Q;�0���n;��F�쵎���u^��LY�rN��t"O]�t��m�U��,���g��U-�eR"DS�9�!|�$�Z)0�>���.�$4��Ŗ��3�ht
��W�$:�-�Vb� ��.��y7�N&�z�0!���
���U�2�gŜn��gņ��nךSi/[��"��?u�F��%��>�g��U-�e��?���s��ʟ0BSuQYy]V$'��d��l~uQ��)���
�z�}
m����TԒ�@r�ADs�lE��8���/���R���7����X�l�L9P|/��V�P3^�h�c*$�7��d����h���n;��F�쵎���u^��LY�rN��t"O]�t��m%�4AХZ�g��U-�e�?���Fߢ�!|�$��A���q�.�$4��Ŗ��3�ht
��W�$:�-�Vb� ��.��y7�N����5�<&�(u�A:�2�gŜn�]�Ȫ�m�ךSi/[��"��?u�F��%��>�g��U-�e��?���s��ʟ0B$"�@������EtJ�~uQ��)�j��8'C�v
m����TԒ�@r�ADs�lE��8���/���R���7����X�lz+w�] ��KB�O����c*$�7�
��\�� b���n;��F�쵎���u^��LY�rN��t"O]�t��m_�p	z�g��U-�e�����I�!|�$��q�n�t6�.�$4��Ŗ��3�ht
��W�$:�-�Vb� ��.��y7�N>���X],�:���ڕ2�gŜn�TKZ%�)�ךSi/[��"��?u�F��%��>�g��U-�e��?���s��ʟ0B�I�d�9���R��(E~uQ��)��&�:$
m����TԒ�@r�ADs�lE��8���/���R���7����X�l޹$�h���7��~g)(�c*$�7�Md-K V����n;��F�쵎���u^��LY�rN��t"O]�t��mʦ�35S�g��U-�e���5�F���"���u�K�����.�$4��Ŗ��3�ht
��W�$:�-�Vb� ��.��y7�NBH��ȍ�_K����h��2�gŜn�&6ޫ���ךSi/[��"��?u�F��%��>�g��U-�e��?���s��ʟ0B�5��ʨq%g'~V>�ہ~uQ��)�?�I�dl
m����TԒ�@r�ADs�lE��8���/���R���7����X�l_l�?��T�����a�c*$�7����1������n;��F�쵎���u^��LY�rN��t"O]�t��mFf!&���g��U-�eM�c@��{AO7��F�e�6���p'{�\ɬg��sB��ÚTK�}�5/uIT�K�^d��.�$4���A��B��g�T�\ ��PzU|�J�ZQ�����s=��[�n&��6_\W�t!���4�f��[B�.*�� �R�j_�3��4�jm��my$�N��.�$4��Ŗ��3�ht
��W�$:�-�Vb� �[�"R���`��Y���{�jP�k$�)�vxѝ�Ө[]kk�%��V��	��yj�����J`�v�����襰(��Wg�D�a�F=n��f�I��~��^V������_�&3� �iY����öŲ�9C������G�����Hh�7�O[H5�N��{��:>�O�S�r���7�u�����v��o����c
~���r�t)0�u��t�\/^�1�[7.�`lI��>4�vp37Zz�)	��t�i�x��V�n�*��������2�h�(Ӑ߅%�$ԧ{n0n���o�u��@�E{A8iMǓߥ�zI�� �5�Ϡ��)���C�M��(=�Kz[Z#ȥZ�7Q�&`���R���U XR"��gLE�z��XN�Z��hq�����}و,�4�Al��yV���9���
�]�!���~�}�D&�9���
�]�!��	Ǹ�y85��G�P��� � 5����)��d��<Ac�6�o8:4�0fߛn�x���_W�y�#F�Þ�^U{���F���`~Y`���)G�9�ƻ2nua����鍾����ȭG�V���تU�|SI��lMh�5K��T�M�r#�9l$���#G��	�c�4�b���	}�@�}��x\������j,�k�o�r:���o���wu6�kf��!��|�R����f�+�ӊ�_�3U�9f�_T(Z���G7˖��3�ht�A�hYX򬞃o�ϵ&�����t��ݾ-/̤�靤�}ODk��v�A�NF��Ԗ��3�ht	�c�4�b�R�%��{���gZS(m���E�~��?zk��Si��]���gZS(m���E�~��?zk��*���c�	�Ky�F��؈a�������Fu*��^������#*<\/i�\	t�AIU��#��9x��p&�[ǣڬ�,��V�.o)�R���,.��Y(�ѡ恙���.�Y�R���,.�с���Z�|x�5c�@���v�8:��$��� �vL���p�!���Ct�w#��@Ż�&ǥ�̻����.�e�	q�X�Z����D<&9 �����`,9�H�W&��a����3�@[��
�}I�?dX5-��ѓ&��a����3�@[��
�}I�?dW8��N��nj{��z�"�~�¦�Q=�=y w�⽒��Ua�� `�]��[���؈a�����.�� gפ��rA�V�cx�k�×��4m�T�4��r:��
����m��gU����*񏫽�{�{N8!�J�~���i�xh5���h���E`���\�ܢ��,�I<�K��Ԧ���ub�t��I��I������&��ƴ۞���G��k�[ dϠֵ�k���O
S	��~��A�;�LrZ�0m�\����n~�/+?qTY�`�v�����襰(��/��-0v�w�(5��d9`�v�����襰(�����̵��t����m�=�er߮�@�N~��n =�|"�#~� ��X?����Z��N�?�����3�ht�b}���9�����Ψ��Z.Ps_*�GqW�w��fD�ws�nn)0�J	�`%��$�����Z@��o{�K۬Rr����#�̔"v���
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�ħƿ�9c�1��8�h����,����^�V�.�	g�y�gߠ� �`g��q>?�=+��r�1�OG�mA�T��2���-*+�m2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�� �W9���+��l��b�"�݀`A���cbղ%�oCm�Ӵ�@1 T�V	�tL��	f�g���Z����������H�WT�%��D!����ހ��g�R����[����"&�&���VA}�v�a'����\�Z��'�Wa�L��ʻR0�˧���.�E����F�Wy��Drpg�-ΘBdcL�qh�  `C�H��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��6�������1�/��*8�����d�kⲽ��uc7�3��׉󾶓�7��J�����k�*ί��Oi��!�`�(i3x�]�V��!�`�(i3����[5ʞ��Ѵ����������?��)(�"���G����%Ah�%4
>��f���T,�;C@����
;�������kفA-TX�Rj�+s�!���r�mj�1����iRl�CĂ�טx�Kl!Zh��1�4��}�Y�V�v)�	 }��x�y!�`�(i3l0��F��j�ܑ�!@���{]�:94��}=�d��[Ya�<!�`�(i3JHn��z�G�zRT��N���������-#��)�?M��7���E����F�'n�^0o?9+�J���D򭢵�#+����wUP`��dpfV�L��nw�4��P�vzo��f�(�Q*J|�� �`e~���|c����(�a�肢�{l�f|�ό���.Ӳk3�� ?]��i�jZ����R]N�By3��<Z鎬�����V`|��](R�_�';���ͳI�E����F�ҋX����@�ڗe'� ��S
e�CHD�u6�y�J2)V�o��C!T*�q���U�$��	�fѥ�[���В����m8�{� ��S
e�CHD�u6�y�
���t��o��C!T*�q���U�$��	�fѥ�[���В����m8�{� ��S
e�CHD�u6�y�̴K��U��o��C!T*�q���U�$��	�fѥ�[���В����m8�{� ��S
e�CHD�u6�y`�<E�dh�o��C!T*�q���U�$��	�fѥ�[���В����m8�{� ��S
e�CHD�u6�y�=���j�9�o��C!T*�q���U�$��	�fѥ�[���В����m8�{� ��S
e�CHD�u6�y\r���㯄�����
L'���Xw��RN�-#����ێ����F���`�?ӄ'yy��N�iM[zigzA=v)�����5	��]�!��	Ǹ�y85����[��3&��㖏��ś��޾&�\����W�GiGn�بpp��ZG!�*��/qRr��Nb�;�43)�$S.zT4ir�_ː�W�{'e�"�,�>E���TD���rs�i���1L��I�G�C��Y�K�za۬���f��yd�x�2�nR�~1e�������=���
����fbK7͍��|��W&":��s�/���_�~C�8"�5eI�9��&о��#dn�'c�����ze�@yo��K��]�BƠ��q�-��|��ϱ��[��q�{�TD��ό���.ӵ�Q�}�qjZ����R]Yl���#�]�!���=�%���b�ђ��V�(^���TD��ό���.Ӎgt�k�T1d�H�Zc�Yl���#�]�!���\B��V���D��˱�Ui��Q�x�gt�k�T�8?�H���Yl���#�]�!���\B��V���D��˱�Ui��Q�x�gt�k�T�տ�G�9Yl���#�]�!���\B��V���D��˱�Ui��Q�x�gt�k�T�^��	�Yl���#�]�!���\B��V���D��˱�Ui��Q�x�gt�k�T]k�WM��qYl���#�]�!���\B��V���D��˱�Ui��Q�x�gt�k�T��0It�N�By3��<Z鎬����y��|�!�p���!���	��*8�����d�k��q���R�>P�2-i_���F��u=��i:���0��H22�բ��3�������I��'�@�TE�J����Ϸ��$q{�f��a�:&�>��s��%�a���fA���������gb��^ֻ����XP���E�z��6�Y�a��	���~,���஽_`6V�?���VIÙ=�H����볨{x���� ��`A���cbղ%����~���;��������!"�S(�J�ْl��]�B�M:��2�R�)��<|�9�a��!�`�(i37�ܥ��2������\#O���o��z>�n�SSC�	��X�6X���(��O��ɀ"���Q�^�y�����9�!�`�(i3��2A#��a1�z�!�ݢ�u!��+_�i������04Tq�`�����L�+P�X�;Qn�Ix��њuw�@.G5O7� �Bo���+�ހ��g�R�]��-5L�-0���+�A6#�a)*t�\�H_��1��0�WQq~�l)�������5	��]�!��Zˎ�f+� �`e~���|c�����Y������{l�f|�ό���.Ӎ\�H_�����H���J)�lV�����5	��]�!��Zˎ�f+� �`e~�����.Ԭ�(�a�肢�{l�f|�-�`��8�4�%��mz%���=a\��J���� ��S
e�CHD�u6�y�
���t��o��C!T*�q���U�$��	�fѥ�[���В����m8�{�X��R��oC�z�C���K�-)K�7Ê7�E�4'���Xw/���:;aR[�T�.�W���1��k3�� ?9<��WI5�^��	�N�By3��<Z鎬����L�`u�K�˱�Ui��Q�x�\�H_�����H���J�I(ީ��Ųo  ��]�!��k��v�Kp��}�G�@����}_v�P�ڜ;�
_��&�1d�������E��@IE�U��@�ڗe'e�	q�X�Z��`�+N[�;�R������7v����B�X��Q�}�qR� ���{Yl���#�]�!��U(<�i�u3~L�uIş��Y������(�
t�ژq���U�m?��"I��":;�����E��@IE�U��@�ڗe'ג�؁�R�^�d��d}�]2�y�Z鎬����Ĺ#{��/���:;aR[�T�.�W���1��gt�k�T�8?�H���Yl���#�]�!���\B��V���D��˱�Ui��Q�x�&����8�7g�@� :�"B��$I��w��,�,�JL��ބ�W}�Q�p��}�G�@���m?��o=�<*��M�Ǿhm��@IE�U��L$�����/���iP1i���m
��5�(����7���	�%���N�ijU-j�`7G#+��<ͧ�:|[��N�w҅�A�=�8bH���cN�Z�3��b�ђ�3稨�;�<��z��}�
��|�6|�+�� VU+I��X��8����]K�I[K'�/���ד*�hW�w��	�x*�7`��KX�U~�?մ\B�m-�;�?��d�٣�����6>��n���ؕ�)���e��Ʃ:�)�9ό���.�9����T�5eI�9��&���G-��IZ鎬����Y�V��#q����y�^�/m>8Φ��8���ό���.�9����T�5eI�9��&�l�`i�|cZ鎬�����h�l$Nh*��ˁs�W|G�_u�����q�{�]�!���1����m2lk���qɍ�6��I�g�E����FZ鎬����Y�V��#q�9�j^��"I��":;зq8�Ј'���Xwa'�<� \��M��U����	�����+�J��p�VU��J)��� �%��mz%���=a\�N/�蔧ε�ˁs�W|�{4�Y�`>j�5�i ��]�!���\B��V���D��˱�Ui��Q�x��K�Q�2r�"7&��K�-)K��n`5�fK�<ͧ�:|[��N�w҅�A�=�8bH����Q��TF��9�j^��o=�<*��Z.��0�W'���Xw�����C�$��	�fѥ�[���ВZD���zQ��g#���1��u�+�L�)�{�d�٣���,�JL��ބ�W}�Q�p��}�G�@���pzl��a��٪Ō����0It���Q]� _ό���.Ӈ��uj�*&��;�of�Ź�O��)�u����pTOj{��`�mǎ01�E�0�?����'.���t�Li��#g�k����ƃ�D�d���}s��,񥩏��4������]K�I[K'�/���ד*�hW�w��	���F�_"7��٧�\�T�q�>�YŇ=�er߮�R�)��<|�9�a��!�`�(i3�3.�<(�V�B�l�2�����j��j��h@S�@�]_LO!�`�(i3��7A�>�x]��n��G�o�>:��GݔO#�Z/��v
���쨳\�J�n&�������C��������v�Q)��|�jь� �`e~���|c����(�a��N�����WZ1��0�WQ�����8l��k���ڜ;�
_���F�-XX!i�X;p`�� ��S
e���z��P�D�+˨a%�X��R��oC�z�C���"��8�O_s *�XF(R�_�';���ͳI��OO�!�N�� Ќ�e�fK�ࣗf�8T����va�H�9<��WI5.�|Ћz�*�\�H_�����H���J;U�2y���苇��Fe� �`e~��2m����4���;c��Ǫ�X��R��oC�z�C���K�-)K�s *�XF(R�_�'N j�S�,Ĺ�OO�!�N�� Ќ�68�S1`�P�=D�<��va�H�9<��WI5j*�//���C[ g��L(R�_�'��N�i����τ�ͼ���cC�z�C��`���P�C[ g��L(R�_�'�����TD-��ͼ���cC�z�C��}�͙Z%ʒ�$��;�j{���ێ��n=�|-;��f�YɴQ�P�����8$�*�J�2|�Z�F_u-��2)�,���Y�> �������Q�}�qjZ����R]�����ce؏{��ʝ�a�2y�s�wd�ч@�.;�<.�
!I���kb�ALb���s ���/i�q�X��X;p`�d����(NZ�^6ג�؁�R�;#5d���_�I�6�k_O��~E=�IǺ���2j�m��yP4&cY_}�n1�
!I���kR#���V�s ���/i�o=�<*����0:t�u�d����(N2������&����8��I(ީ�����h  �G�at��ʲ���:!�ӊn�&����8�-�a��~OD���K^�)wd�ч@�2tcL����@[�_zβr�v������P�/eոk�j�
��j��Ξ/�H�WY\`��J��-#��)���Q�$��|6�ɚ�!��t�Li��#g�k��{=�RT��Ƙ��}�$��Ml�44]��锴����e���SMI��pA}sJ{=�RT�޶N���$f�=�zD�����锴������h(��"Jk�\�)���:�ߧ�������R�����-���(u������ m6Vhj�;\E���'#@���q�ڜy_*t5~p��v�w���WUI[��-���(�=`�x%�gt�k�TX�����P�`�?ӄ'yyl��WC({=�RT�ޫ��K#i�\���	��6�pl$�1V��	��yD��+?oB{=�RT����OL�������9C������' !ǥk�}���v�i'ܮ�f$�(l��{�ot���^���\�}5eI�9��&������%!����ل�yx��}� ���{�8	lc�*of5eI�9��&PͶ�����\,���p�����ل��8��V\�ƘZ��<5�T����_�*(� 0�p}��4ܧ1`�?ӄ'yy~��y�\�7����{��=a�F�Aߥ6����b�ђ���)�r���O��8@�����0�wd�ч@�l0K�VWe���Ni����8�V��a*��4�磕5eI�9��&l}
@Ŧ`�?ӄ'yy��s��nM*)��g>�����s���	 X��-���Rv��\�F\��D$�]TF�F�������8���^�蚍�6��I�g��`|��%kr$(��_�2r�"7&�a�
��5���1��u��P�e�jXҴ���G��2�n�Õ�&o=�<*�ւS���FO]�b��ގ�q�~�Jf�0h�5e�n`�@b/ἓ���h�ѱ�����@/��r ��H�7�%r�ϱ��[���(@CPw5eI�9��&�\����l��Q�}�qjZ����R]�<�t�yx��}� ����<���b�ђ؏�` t�:�5eI�9��&#����[��gt�k�T1d�H�Zc��q9+t�}8$�*�J�O��~E=�I�jʱ?��s��ɛ�?өd����(N�1����c�Z�~�&����8�Lc�Ո�D2��$�\%e���<���k��0:�3ә&�M�4�Mv!���x��˓#����:��0^�d��d}_?��Ӛ�NÄ.dW8$�*�J���6��I�g�S����&��tv�Ҹ�z��ic�ג�؁�R��"��8�O__?��Ӛ�m5�8$�*�J��s0P_!�S����
�Vw�*��ᱪuuג�؁�R�;#5d���_?��Ӛ5��ܴ>���<泩���;//��` t�:��2r�"7&��H�ͺY���gt�k�T�^��	����	ΰ�A�.�p��N�J�d����(N���<&h�:��6���I(ީ���𭨈��� 4�04�jf��ܐ�}ļ?E�!$6ӊ��{��t��MJT�G�荸���th�t�X.S���������6tMk�j�j#��t��MJT�s��0X�wb2�Q��Q;�im��ɝ\�!2A�߻ ��Ǵ=��d%�Z9!�`�(i3���)�>��hbV�֎c�(�.�����5f�, 쪺.C�`:��Q1e���ZYM	���`6��[(�4���/��NO�l����m�=�er߮�P`��dpfV�L��nw�4��P�vzo��f�(��q��P��X��R��o�J�"9���^�d��d}s *�XF(R�_�'2|�Z�F_u��OO�!�N�� Ќ�ΰ��$<�Ӥ��,V����va�H�]��i텅ir����\�H_�����H���J)�lV�苇��Fe� �`e~�����.���G�t��� ��S
e�CHD�u6�y�J2)V�&��^wڜ;�
_�ʇ0Z����C[ g��L(R�_�'O��~E=�Iu�$��-vͼ���cC�z�C��t���Q��D�\�H_�����H���J7g�@� :�苇��Fe� �`e~���F�TY�~ox�t�� ��S
e�CHD�u6�y`�<E�dh�&��^wڜ;�
_��o=�<*��QY�\H9�� �`e~��2m����4�+�L�)�{N�����WZ���H���J�I(ީ��ŭ`'�n�>o� �`e~�����.�����KD4N�����WZ���H���J1���:[�o� �U�O��/�g�W�G,�?������7����yퟻ T�٪+_3~L�uIŬ�(�a��(Kԙ+�΢#�$���8$�*�J���6��I�g-��ȴ��{�څir�����&����8�)�lV�k��r�
�Vw�{Ē���ג�؁�R�^�d��d}�,����N}��a�_���Xj^6�	at��ʲ���ȍ�)0f�(Kԙ+�΢5��ܴ>�t��)��^����;//�[���U?�]~� M=R#���V�s ���/i�o=�<*����0:t�u��2r�"7&����^rg��s ���/i�]�b��ގ`ڱR̒�2r�"7&�`���P�8$�*�J������TD-���٪Ō��&�$,��8qTmI(x;��|B"�޾8����C�u�RvR�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯�^��N�&��?�2�1p���}������]�0�lK'���Xw��_
�u��>Oʉ��R���=ە���oH��O>�Y�<]/2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���[�}c��G+�
�c�~9�[vĄ4Ȝ"nF^�_[� h��.c��^�
E�;�#�%�R�J9S� �bRw�����IL�+��V+Ƨ�
}	��Rk�Q[��0�_��F�Ll44`�D�dl~�E���9�PJ���9�ׇӭ��!�`�(i3f���Ն�t�P҃�G����f8�C�XS�6��VA}�v�a'����\�Z��'�Wa�L��ʻR0�˧���.�E����F�Wy��Drpg�-ΘBdcL�qh�  `C�H��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��6�������1�/��*8�����d�k��V}�sw-C6%K�pı�6G2�`e�V�s#��ْl��]�B����=���hbV�֎c�(#nk��"�,�>E��4];ˍH�!�`�(i3��:L��:���H������5f�, 쪺.C�`:��Q1l0��F��jY_���P[V����(�"����W
	6K��?r	�'3��s��'l�X�~g�3�Р���A��(!1�9�͆�i�����%0� ��ۛS�*H���	��<�����`�+N��B0�J�
�:�I��&��)�؊��i�1aڜ;�
_��j�;\E���Y%T��BPS�)37J*u��l�M�Ϥ �`e~���|c�����Y������{l�f|�ό���.Ӳk3�� ?9<��WI5�1!u7}:N�By3��<Z鎬�����V`|��](R�_�'�s0P_!�E����F�ҋX����|P�������A�=�8bH��&��ѿ9�(R�_�'O��~E=�I�t�5ńҋX����|P�������A�=�8bH��&��ѿ9�(R�_�'N j�S�,��E����F�ҋX����|P�������A�=�8bH��&��ѿ9�(R�_�'��A�.�p ��H�Q�ҋX����|P�������A�=�8bH��&��ѿ9�(R�_�'��N�ijU-j�`�ҋX����|P�������A�=�8bH��&��ѿ9�(R�_�'�����TD�E����F7G#+��Q2�+�Y�{�rN�cZ����d�k��v�N��!��`A���+@�����_�>+�J2)V�����
L'���Xwo+
�B���F�-XX!i�����E��@IE�U��@�ڗe'd����(Ns�yze�Zv�����
L'���Xwo+
�B��q�X������E��@IE�U��|P�������A�=�8bH��&��9��hUO��~E=�I�t�5�7G#+������z����A�b�*܋����V	2M3����;//�V�(^���TD��-�`��8�4�%��mz%���=a\�S����=�����^�bp��RP=	P��(�
t�ژq���U�$��	�fѥ�[���В����m8�{d����(N�=���j�9�����
L'���Xw/���:;aR[�T�.�W���1�ג�؁�R�^�j���7Ê7�E�4'���XwI<��f�?��6�J=�A��Y纽����8no^�#ҫzU�	vn���-U%�o����, ��� Oag�qod�֓���`A���cbղ%����~���;��������!"5�d#.��?T�]D�9�"��0��t�_[�v���U(�M�z�ۍ�1k�
��o��C!T*�q���U�J�"+?�e������]�!��.^�@CGH9M\��e2��p-!]�5y�����胬<ċI�wb�H��J2)V���+�J���q���U�pzl��a���gE���؏{��ʝ΁�a�n���n`5�fK�Q2�+�Y�kѶ���� k���3"I��":;!�`�(i3�d�٣�����6>����9וP�;xB�_/1d�H�Zc��E����FZ鎬����Y�V��#q胬<ċIX3�A���\�̴K��Uֲ��+�J���q���U�pzl��a���gE�����JԶ�.�$#e���:�n`5�fK�Q2�+�Y�kѶ���� k���3]�b��ގ���V����d�٣�����6>��؇g��,�I���$D3�f^�E����FZ鎬����Y�V��#q��]��A�k���3�z�Q�q���+�J���q���U�pzl��a���N�)�-�;�Eo��K��]�q��n`5�fK�Q2�+�Y�K=J��(��oM{r!:�k���3�z�Q�q�d�٣�����6>��P��r��c�y/=v����;�Eo��K.�wK��� Z鎬����Y�V��#q��d�M>U9��
�;�Eo��K�C�p2O�q���U�pzl��a�D���"��	���,��bJ�e�C��w��z䮃��Qi��+���>^�#`����V�a��6G1��xY?�B�l�2�ՉSu'�#K~%+n�=�ͥd��7�׍���ebCb���]3�1P'��:DE��Z�h]�3����k�*�q>��`�j��5��o�	P��o%z5��ܴ>���o�32/�;|��T;�v�$���;Aٮ!�\����qjI~���ʳ���GJii�"_�`��-:���h�@nJ���t�#TV�� x=3���R�V5j�Ć�O%r=��E�]\�
�Q�}!Z�Ő6?#�h����(J�F���֦VE���T�8���p�l��@��5�S�5��ܴ>��z����Pڜ;�
_��5��ܴ>�:�}��E5��i�7�^�f`�3�y���n���>���ɑ4Y��u�	"Ocbղ%�R��GN@����x�hn�B�l�2�����^t+�
�<ݬ�KfHړ׼[QR�)��<|+!N�e[�������"&��2�U;��|BtZV#�z~j�;\E���!�`�(i3W��J�}1��0�WQv���?����Q�}�qjZ����R]����;qͼ���c�J�"9����d��Kd����(Ns�yze�Zv�qr�~�룤 �`e~�����.��U"Y+р�M�����(@CPw� ��S
e�CHD�u6�y�y�8�A�m��yP4&w�������ͼ���cC�z�C���H�ͺY��d����(N|u��W�s���6+9<��WI5Z^ >�jPF]�J��I(ީ���:��͟4�(R�_�'��N�i�wK��&6j�"Hs��Scy!9x�����A��Y纽&8��U�W�gSS�[nl,m��#���Sg�W[�E���j�,+$\�M��lJY�Pt�-9VFg����R�?d������X.S�����W�����C�"��0�����k�*�.�a�n'��@	J�!�WW�+���3��0��A����}������"&��2�U;��|B��w\�'L�O�*]@!Q$)֫��)B�	�>�D�J..�E���?��)(�"�ސE}yޱ;��|Bn��[�2|�Z�F_u!�`�(i3{�R�$�Vք ��S
e���z��P�*��ᱪuu��_�>+�Sծ��[�$�
!O:0��kU����Y1��0�WQ�Y'#4���&����8�)�lVJ�a$�Y M�XtM�N�� Ќ�z���O���t.�M��b�ђ؏�` t�:�;?%���ڜ;�
_���m5�m?��q�X��N���&U2�0�FOQPg9<��WI51X�����gt�k�T�տ�G�9{�R�$�Vք ��S
e�CHD�u6�y��`���d����(N|u��W�sM�XtM�N�� Ќ�68�S1`t��+�}�d����(N���<&hM�XtM�N�� Ќ�5M�N�]�o`o���կ�����,�ǰ	M,��rERO�*]@!Q$)֫��)B�ߘk��-o����І=�ra6yD�� ��p[�ٕ����se�{�z��x� ]
�<�2�Ҧ1���Z�וN�!��-�:G�]�����<�6^١�Z�D2���w`�����.^����"�~�Y,�9���uS�����@���\�dU��Xp���ڛ|J�PъT紒�)%��ݼ�y�:9�9��;�x��������0�e��6ڿ ���M�M]?��f���r 	�1���/S|Lue��Yz���A��1q$7�#�Qk�v����<4C_����n�[��*�H`�~�ܝ	�@���oR��5l��5���S���\NG�1dɑ����a�Vy��LAF�����nĠ#��t21Fp4���Y-��+�=S�vʐ̿y�P��8��6���|�;;�
�����0�����^B����Ыl���#%a`Y��GU��|��sk/ ���ѡ�*�|lC�y�ZDU�.��%��	����D����_�̈́V����?��Q/�����3�=�Z�����r
 �;)���x����Y��Zn~�EK�l�t.ɣ���z
-��|o��f��wN�$z��+��o�u�/���g(��
k����:�F7��3볒��-���6�J��ʒ��қ{`Y��GU�X`��_/�O'{��In��2�8.�xy��)�\�1�����r�9�>���y��&�/|h&jquP�������L<2<����*�|lC�y�ZDU�.�S�<���壦Zw��!�nٚ�2�,��qi�C��U�����C�w��o�GMG�2�3�yc�A�̍�)�y�YWYdU��Xp���ڛ|Jľv�鳔��3)$�f*��T%������yC��r�sl���o�u�/�1V*���p�mf�{��l\6�he�o"x�ȥ�i'�˳�ݏ1����:�I��&E��-��q��H}B�úY�t5���̔���;�77:�2��ɉ���Mβ�^�/���-n�9�U~�E)�GJ�G#����Z[��<�z�qT��m��zP���	Oe�ُ�AH��tnZ	�ɬb�H/��G!�����3�i�r�Թ
5�ϱ��[���(@CPw;?%���ڜ;�
_�ʯNÄ.dW@�uU� �ꖱ_�5���M�Մ���"�,ݤ �`e~���|c��/)����[k���3"I��":;�N���&U2�0�FOQPg9<��WI5�6�昆�r45�`�����(�v.2`<���/Է0c(���(R�_�'�s0P_!�3���?�xB�_/�տ�G�9{�R�$�Vք ��S
e�CHD�u6�y��`���И|��,��A�.�p��ּkU����Y���H���JLc�Ո�D2�3���?�xB�_/]k�WM��q{�R�$�Vք ��S
e�CHD�u6�y����ȫ_V�d^_�Rꑽ,�I�t:��h����b�y��־�U��sp֟kh�W�f����C;��҇И|��,2|�Z�F_u��â��E�❽�J!�z*�9㞬|�M��5�М�\C�)1�ﻙ':]J�y�ZDU�.��2��[�rR�Z3�@�GݔO#�Z/��v
���M�wScp�)Z����(k���3���"�_�iPL�@�tj�(��d.��H�f�ȥ,�rXK-�?~�S��G���/�>RT�>'W����Ŵy����O�!7y�x�}�0�.�,�C��A��L��޹��LU�L���b�ALb�����}��a�G����)i�,�I�R=]�}8a!n�}'n����wt��j^E�z�G��1vo��W�y����O�!7y�x�}�0�.�,�C��A��L��޹��LU�L�������T'.��}��a�G��_��M� v?b���7;�Eo��K�>�0�З)0kcj1�kD�������r�y����O�!7y�x�}�0�.�,�C��A��L��޹��LU�L���R#���V���}��a�G��_��M�y/=v����;�Eo��K�p��h׬V�!+���}9��m;�nJc�='�k�rR�Z3�@�GݔO#�Z/��v
���M�wScp�)Z����(k���3o=�<*�� �������c%����o=�<*���!��4@ȥ,�rXK-�?~�S��G���/�>RT�>'W���y�l��N�PΚ��_�(f���i�t�U�<�S7���6I��|O/xB�_/]k�WM��q��â��E���h�e�I(ީ���a41h��ȥ,�rXK-�?~�S���Q�}�qR� ���{w?�W�S[И|��,"��7Ch�m��Q�}�qjZ����R]xAp��4 И|��,"��7Ch�m�gt�k�T�1!u7}:��>�!觪И|��,"��7Ch�m�gt�k�T1d�H�Zc� U�����pZ�pF�l�J�e�C�ꞼV��;�G�����;//��` t�:�yg��c|q!И|��,"��7Ch�m�gt�k�T�^��	� U�����p�T��i�LU�L�����ج�~|�d����(N���<&hy75���ri����a�9�;�Eo��K9=�-���EV��	��y ��f"����A��(aMq�P���p��/�4�X�q�	��؄�e��c�쪺.C֡�mG�[�}M��0�d(_\�^?'qKy���\N}zp�jN�^�_�~]x_/�Z�s:��T�����E�ȴ�TΉ�6Rρ\=ʺ"���c�
+,I�20a���ac������,!��?d������X.S������}q����:'��HV|��V�a ���Ɋ�ZS�[*�$��f�z���H@�{�'IK�L�����d�kⲭ��2F���3��0���wȝ�G �VL�(\F2#���h�黩~�S���3��0���wȝ�Gھ\f;vM�*��ъ?�i�;�>�fͅ�ݮ��a�=��d%�Z9����r����<���黩~�S���3��0���wȝ�G"�����'��]a��z��黩~�S���3��0���wȝ�G"�����'�z�	���黩~�S���3��0���wȝ�Gھ\f;vM�㚄��ɌTY��G�Ie�i�(R�_�'�����TD��W_�`��aH�J H\�@[�_zβrB�ek�5W��ɑ4Y��u�	"O��3R~r��&8��U�W�gSS�[nl,m��#�Q�%Z��;&�����O�h��~x�۶�kvɻ[?�V��!9x�����c6�c��A>	�x��FR��GN@����x�hn�B�l�2�T���)� �r�hr�W��xO@��U��ݮ��a�=��d%�Z9ھ\f;vM�*��ъ?�������H�ݮ��a�=��d%�Z9 �VL�(\<e_XP�v1��ԏ��R�)��<|k�݈�x�L�:��aqV��S�Q�z�
߉�T&8�hbV�֎c�k�q��l�czD�k�$8�2�-Me���qfb�B�l�2�e�St�F��6��ޡ+W�9u`�w��UAV�?�� �`e~�����.�uK[~�H�įԫ���\�g:Ļ����,�ǰ�M��%�$���%Ὠ�p���\���`�+N������@n��C��ip