��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�Jз&�6��`�,�2����yׁ @'�إ��(�q�<������0T-~�	�Y\�������/�'o��Ӻ��,Q�Q�?uG�Qy����JN�YQ���b`.�]2'%Sǘ+�����I�'�z��9���
cC��O�-��G�s���R����#1X�.ՅT��+Ϩ1Q�2�:C�.0q1��B�ce�jͻ��}�����9�Kو��. z��ڠ�1p�W��b࢞�i�Ot���k`��$r�^�A%�7��� ��R�āy����yoZ�P/b^��GAjc*!�� �]K�lh��.��:H�T�fޮ��Ĉ;��~h��h�W��>�:��)�򹉓��#�)��#�)�� A�}Z�n��-�4�E͉�-�DfWn~��7��+�gE��e��d*��N���9׬��Lw�E*��+.3����sv�RS�6�1M���yK����ॶE*��+.�}���n9��W�Mށtd؈��k�;4���Fz�	�$C�jQT	�$C�jQT��x���t���R=l�#�	�����g�Έ坩� <�44��v��,X���.�bI	\����	d�ዊ}��~:�u���n9��W>X[V��k"Y��^4~B+�9�'���Fz���Fj���Fj���x���ti�8P�-�׭{6V_��J&���1�c�ؒ,�X���2���O�hf>Ŋ�g��@���"�Q�8t�s�0���8��t�\����1�x���0��%C��0̉YaA�=̮Bq���'�y䜠�:�A�}_�r�t#�+��O��oy��09�nXm:m�t
�W_���1�o��Sl�xdG�!�5��� ��YY_���6�z�
^��1���K���π�>���cl8)��� ��J��b2�K\��$����\O%���F{�? ��:��c�b����f��Y�5�7cWr��
�1�ِ�E㟪g�7�������0A�OT<��y���@��v�m�qs,�Y[Ն�l��"F6 崭��oes���$q��mKx"E&��� �$Y��C��s7Ҹ���/JF[B����,q�.3��h�V�*�U<������P�S�bN��4( �.x�����fg��ͥ������QH�<�h�d���@빮��1o���W+N��<�DU]sȸ�"rR!�`�(i3VR��|B���D���
�չ	L~�BA�kN��&94$2�¤}l����Fvf����P��~w����+���m@�p�Y:
�B'���a(G����h+=o���&>�S�䡢��k͝�ul���C�A:���i�����Fz�!�`�(i3��^�j��VR��|B���D���
�չ	L~�BA�kN��&94$2�¤}l����Fv+�-EP,]�!�`�(i3������=O�Z�:���ro�؛�36�ZpMu�IRIn����\'tI�D��ܛ	g�p}XR6��^U���Y!�W�Vc�sNL�u�
��Xx����G�$�-7좎E&(p�
����d�k�ViR��W�ik2)�
}wʭU&H�1��8�h7H�u�ÍeZ8��
;��d��q�G�a�P;m̳�UlgRQ�t|Y�f�sJ�F���s�V�����<o�nïi�JHn��z��r9�3,�qo�,ܛ�	��|��	(���zL͊�q���b�Kzb�d&(C�#�7#^�Vn�^ֻ����XP�����-����[�f;q�sɈf�=K����X���`>;�`w��^e@��V��M�P�zL͊�q��o���.N�wJ�G�����t �JHn��z�w٩L7���i�^e	�F�K����'�Z������be�o
85�C`+�9���m@�p����
��s6��\�v��wc�}�![W ��"vY0Jߺ�'n�^0o��]�mj:�ǆ�0��n-=1�BF�k͝���<���r�����z5Ā�����^�j��C �H?�o�ݷ�����.j�,�3*������|���kJ�|��].��'���Xw����l���(���e���!n}y��Y�{'%s��.|Z�����@	Q^�V]��}R�wX��*��p��U�d�K��@�!n}y��Y�{'%s43u�R��}/A;T�c���Y#?M��^e@��V�m�C��x�T�\ ��fȂ?�x0�C�Z���8k>6s����]�!��$��lW�d&��b8��)R�v�w\�L~΄gO�3f��*����f���,�LoG�ٳ��?T�]D�9�ϑ��[��;e7�)norǟD�uiL${?�����>��yܛ�	��|��	(���zL͊�q���19TH���'�3�$ �#^�Vn�^ֻ����XP��Ȼ4�t=�j�.�/'�����W;5B5Y+� �i7�sp>�O����!;�Y"f��g�o&�Y��>�_���ˍW�}�ke�Ts
��q{�f��a�/������#��=ό������?*	�ML�벗0�HC�a*�u�&� LK�a�]G��wi�bZ��b�Bv�~������]�!��%��rSe�u�heJ��Dv�~������]�!��ߌ�>!�0ӆu�۲.��!n}y���q���U��@���Ϧ��Ig`i�ҋX����@�ڗe'�D��/���_3#ڸZ鎬����R;j?�鴜�֞W��{l�f|�ό���.�c�{dϨ��B�>�9�6�vg;Je'���Xw>\��p}�	��D܂�A݁ؠː� ^��y�C�9a<�YVKsz�D�W��Bc�i}3�J��؈��k�;4��K�Q8@"��_o�'�Sx�lޞ��rs�i�jf� l�ǉ��F1x,0=]^	�&������$Y��C��|4�ȟ�|Q�P���2��d�٣��c�A�L'��!�a�&H�[&-n�g��U-�e5��e6²W����_]g��
F�UTz�`�J�'���Xw�j�7����ӳ�Y�
X��������`y���pzl��a���#�NN�y�����Ӑﻋ-�����S8�/ #O�)��BT�^��a(􆿳���L��F[q磫��<�:�π&KXҷ�YdS�=��6��+ͻ#q�H!l�5w"^	����3�K���蜍6���Mf���9��Y�{'%s��.|Z�����@	Q^�V]��}R�wX����K�Q�LP.���.�D�m �Oh��M�aQ�q���U�pzl��a�&W4�b�A�w���, n}]�}��V'���Xwa'�<� \��5"�7t�J�4Is*�I94�0.��=Y��_�0z�cUL�%*��"����A|��`y����s��d�\��MN����!I/�������A��X�@�5��6�l��s�����[� y�~��ż3���F����T�O�H'�J�����=<�HI����>�W�_=��0���̏�u�=Cm�v4��61��7a	�����Y�
ɸ�oƴd��t�'��9ܛ�	���V[�+
�l掝�K\m��U}�	|^�׽R�s�DH}�_z�9�E�\����8�i�`!31u{w�S� H"�nT��z��uWU4y5=>F/ġ"���Չ-RW!�՗"$p\�>���S�w҄�^��(I�>'����	4T���\�nƨP�ʱ:��Ԩ�\�"ߗtl%�]Y�%���Ádo�d�x��u�5�h�br���lpda���?̕U�/j�g4A���{0Yafk��r.y����nL���~C�V�T��a׈Eg#f�z�q���<�{�!���"4��:@��o���KEd��]^X0��
x-	���'�$HgL��)������e��Q�Q&I`��=J'����r
���I}}3M�C,����|#^�Vn��l�M�c���=^��>D�c�lQ�����+�7끍J�[T�)��o�B��^�֌���<�a)�m�d�so�}a�C�ub;�;���dMb3���y�z�ۼ��uWU4y5=>F/ġ"���Չ-RW!�՗"$p\�>���S�w҄����vd������	4T���\�nƨP�ʱ:��ԝ�XLVt����G��5�&��p���P�#�|�B�X�g�i0\��.�gIt�!�����o����x�ҡ-�ّ�^ $� 'fa�#�i~0!�r�qU���Qv�EoO�؁'/B{�;4fx��V$�w�}MX�]y�y�3�˝��28Zlۨ�\�"ߗt$��6�iy��7I��XG��]�w9"x�g�Hz���MN����!I/�������A��1��+�W�Ń�I��-Nd�����R��Y�4��'�i��؏��]�R}BK�ߋ,D���@�wR�� ������tY���F���ø��$�&$�^��$f8���]�5]~^�����L}c��my����d|di};�_͠E:\��R��-=D�`��X~wU2K� ��uF��	Z�����i�r�?�y)��0�0�h��#g�k��G��⃵V���A=�aY��m[�c�Z�~�]X����Ǵݵ��9K;�-~i��؏��7��gRv"@ыQ�\b �`MoqF}.	�jo���wJ�G�����|�q<�_��s�֙f�P_�<�ey;���W�b�aY��m[�=�<�^����,�ǰ.^�L�q��D���K�����ƀAh���b��hN8���U���-�?,��/T}��]�?�y)��0�0�h��#g�k��"����J�=O���[�_7��ҩ���xsq��?�d���&�X�'�(+,:ZG�;�d�]7��gRv"@��/��rS�#�g�\&A(`#{��0�ĸ�ٴ֍	��Z:o��|��2��O\���|F3b��ŲNGl�(�	�n)&=O���[����	_ȥ*�sk�NUc�C>���ӳ�Y�
��m_�\��MM
��,={H�3)-�Q�H�����p��2d]o
��?�4b"����~[r�&�mر�R'@�D�x�:�gңs�K�2AYc��V��$���Y#�5[u��Ƴ��^e@��V	g���w��T�\�@��ѥ�+Ȑ�b� P:��s��a�aj�E�>��wL��4�̍%��v�� �F�F�$L���������"�׼L:�%��9�]�3����s�]�<ܥ��QEU����@�LP.���.�D�m �Oh�����9#�����Y���S�@�v��z�(Ԭ�����`^�	�S�_���k�:|�P��� �F�F�$LF�!��T%̵P�B-�\&A(`#����c�Z�ٹ!5�j�BEޥ�8{��$����E`���Fi��|�3;c�<��BY�B�0󕹎@�m�$�b@a)�rg��	8��3�1��y��I{GKg%�+J��nX:F3�s8��q
���E��	_H�#�4�8��0�uu+��Fz��pC��)Va.�e�H�5�	����{�)`_46C���n�SU��\5�OYp� A��!A�cU���?*��|����'3�J~��k���)ga��<ta0������]+���w�f�:�#Wҏ�`�+��b���ف�<5�NlA�c������
��Όú}�s��K j?4��6r_�a��	��$?�c	�| �ɭby��aOw�#�S�&ʺ/�蟞w��g�+�Ĳ�6wK���,���@عE^��8�ޕh�X�7�ЋD��R#c�!��.ЌY�ߓF��A���8D�K^o�B�
/Sq�r��2#�
��/�;�f����@	Q��[�Fc�k��˚����Z��c��~U��|KG?�8&�Ms����g��������k�<DC����?�B�I:׷�F׫�J��l� �[��׍����������*���3m��U}�	�2�G�Ml\P�O����X�e�6<�AT];@���U@���:��F���Ed8���d&(C�#�7#^�Vn�uQl��wJ�G�����t ��,������?�y)��ww��{"]�/ښ[T�r Ъ��ا����20q� \��l�(f���/Ax��}*����>zO�bZ��b�Be��ڡ7o�u��Ö�]���ƻ��q&�<ν$�[���Έ���� ���ۧc��YfT &�t�uÓ�h;���mFw k�1���=���ۧc���OV�ԼNo�uÓ�h;	��3�f����vV�㉨���(���%h���O�v��
F�U����͏ޭ�\������h4c�LU46�����z�C�o.t '����X�*N/�p��<�*�n���wFH���}��a\�����锴�;��|B���	��+?�d���&�O�ʬ�'�~'�f�H�0��̌��"� #�g{uI���l��1��9ЌY�ߓF�ض�g�o��<���g<�\^���\�}L��faNV�T�[��6���ӳ�Y�
��m_�\��MM
��,=?�d���&���e#��2�T�MJ� L[Cv�h�x�l��1/Ax��}*� ��i�cY�7a	��������W5�\tCՌV�����,����_q�_���13�[T�)���V��ÑR K�R����Uܛ�	���G�˹Ď�r�^K������О.�����@���U@���:��F�6<�AT];�q9�+_���	��f�\��=ښ�P�S�bN�CS��ejl�;�w���h���X �d9{U�p�W�Px:'0c�jv�Тk�=�er߮�+�zN����!��ZB��M��7A���:ku��ՁO�#dh���X ��GR�D^p�U�����8M]x�h�h���X �8@"���ⵛ���p�U�����(��h���X �8@"���Y?7����ۧc����D�d�[r�uÓ�h;������k�?�N�㉨���6��0���O�v�0�V��V�2��-�F�ܴd��I hZ଻|��{�Ln���WN�d7B�����P��g�V��	��y�wK��&6j�"Hs��S�<뒯�,2�&8�uP�T�U:Ϛj-��8Ljgޠ.�5�Ϡ��)����jJ����O�n5�\�3��QMWB���t���tH����������P&�wf�3 �٩\�YЌY�ߓF��A���8D�K^oO�[�]�����n*1�#�;�w`f�<86̣��t���/��=-�� �F���n��뾦�6�`���V�#�-K���Ӊ��F1x
�ߴm�>�C�;��_�t��s����?��;��W�X��-��4�n
V~$�����lJ�4Is*�(�����!�+���8�׏�����M�(�V�ܼ���s��߸��S�Ȍq�n��	3�J~��k+t���تa*]R��������56j�"Hs��S�<뒯�]OF��K����0�=��V��������K��S��Q'��t|<�kf�:ҹ���7��q���8���^�d�}|c�q{�:�¸��o6x��i0yXr#�9l$�5[�M��8�|����xP�Q����!��|c�q{�:���k	��F/s}�]�����
��RR�,UO��Ⱥ��#��]��C�1��"�J���Ę��(h�2��}/\�^&%≉=���ʞRػ�[�會1@��
�2`�֔A1٦�+�m�`�+GUz��n|a$E�k����N�V�wvp�T�$3]]��?"|�q�r��<�����]�~�\e����w�X�a���>���`����������n��脯?k~�CV�M�·zB�dR?lPku�O�f Kt��QctIo���C�� TḾK��B�jC�T�٩\�YЌY�ߓF�ض�g�o��<���g<�\^���\�}+���Ã��n�&�E�2�_����0h�5e�iԄgc5E.E@�Z'�^����	�c�4�b���fΌ;i���@	Q��[�Fc�k9���.:���؈a������]x{^���wFH�����b�n�yX��WG ��o�J��p�a*]R���ZHOh#�ï�ɛ�?ө�5ߧE4��
��T���x�;	㯰�$�)�vx�(�W��S#/��=-����7;�gw-[X-���$V���Z�%�΁�Y�<	�����+���Ãp8,3s"B� ��~��	�c�4�b�l�;�w�����g�������5m��l�;�w���d)��X]c_�t��s��1B"�A�`�=�ȭ^0E���^��0�$�ð��Ts䐼�D��4���f�	��kU5�}��N��]���/D�iԄgc5E.E@�Z3F�c���W�x+Q�**|���.�Mg.6�k�5ߧE4��
��T���x�;	㯰�$�)�vxc/���[��WN�d7$V���Z�%�΁�Y�ה��+���F@�m`"F�}�y��Ps_*�Gq�p���x"��`�Z�SQ4O�D�-���f�euq����"���-��$�\X�+Qo��ʺR8���ҳ�N�F�-:���h���=<�HI�^j�iʄ�Ү���<MzD�M>b�B�2����y��l��%����C�Uuh���#� �Vj����C$/U9��H�+�[�q��&d��_2G��T�!����ԄUq �'�{2D{��E�g�@mLq=��-�ju�����cC�	mp)̐뢓e�L;VGdd)ʃ�������?GQ�.��V��?oj0V5����'�u�W9PN�@B�{!d�����~����p5��B�&�p �᠀P�����i��ӯ�0�<��A/%�V�>E %�1��(��2Ǌ>Jv�F�����u�t����-��z
�E'����s�d�(����{�QF���.v�F�����u�t����-��z� ���ǒ,���s�d�(����{�~��P}Fj*v�F�����u�t����-��z���P *���s�d�(����{��1M���yK,΅kit�ϋ�4�L)�ll�X[R��Μ�٣1�"���i�My����G���C��V�RDFR7�EH`�1�&�(���̠�(�B�'`�J���x�����S�Ql`2��~�]r����#�����=%}������G�ۄ��O���azhݪm����Y�{'%s��c2]�l��aC�h�>3�@d �v��t=��,\ަ�Itu�h�ɟ�B�I:׷�F׫�J��q{�f��a�:&�>��s���� T�8m��U}�	KݗZ:���'n�^0o����y�]@���U@���:��F���V!���IÙ=�H�����h<����m@�p����
��s6��\�vūx`��:�W ��"vY0Jߺ�'n�^0o��]�mj:�ǆ�0��n-=1�BF�k͝�w �I��!�udݸn�Ѡ�i�L샾�Q�0�	�A�����<��z��}�Q2�+�Y���awf���Ig`i�ҋX����@�ڗe'ņA2c�`��|��].��'���Xw��*9����Ig`i�ҋX����@�ڗe'�D�6-�˄�|��].��'���Xw�s����5��Ig`i�ҋX����@�ڗe'g��?`-ʂE�����7G#+���[H��8U#��L��G��l`��q�P ڨ��S���Q�V�ɶ�w��I�����q�@��C����~ ��=�F�nܰ
e"��Y�č�Y���S�)37J*u�38BqN�S�E��l���Ig`i�ҋX�������!S^d�z��,�Č��M�x�q���U�>�����w̸���ǃ��|��].��'���Xwk���Rs�f{ �$���{l�f|�ό���.ӦeC���^A e8�~����(�
t��p�VU��J|�+�� VU+I���htf�g�	F�1!��̩<�){:��=Y��_Q2�+�Y�$Y��C�?}�V��Y��=Y��_Q2�+�Y�$Y��C멱c�n��y��=Y��_Q2�+�Y�}ϼ 8���灊� OgD���g9Z鎬����Y�V��#qi&oKo�3r����=Y��_Q2�+�Y�K=J��(��,����NSx�lޞ�ό���.���K�Q��ƹ���hx���X�d�٣�����6>����<2 ��N��WN�d7[B�����'���Xwa'�<� \`h6]G�����x��d�٣�����6>����&r!ť�WN�d7[B�����'���Xw�6%j_�z��MN����!I/�������A��X�@�5��6�l��s�����[� y�~��ż3���F����T�O�H'�J�����=<�HI����>�W�_=��0���̏�u�=Cm�v4��61��7a	�����Y�
ɸ�oƴd��t�'��9ܛ�	���V[�+
�l掝�K\m��U}�	|^�׽R�s�DH}�_z�9�E�\����8�i�`!31u{w�S� H"�nT��z��uWU4y5=>F/ġ"���Չ-RW!�՗"$p\�>���S�w҄�^��(I�>'����	4T���\�nƨP�ʱ:��Ԩ�\�"ߗtl%�]Y�%���Ádo�d�x��u�5�h�br���lpda���?̕U�/j�g4A���{0Yafk��r.y����nL���~C�V�T��a׈Eg#f�z�q���<�{�!���"4��:@��o���KEd��]^X0��
x-	���'�$HgL��)������e��Q�Q&I`��=J'����r
���I}}3M�C,����|#^�Vn��l�M�c���=^��>D�c�lQ�����+�7끍J�[T�)��o�B��^�֌���<�a)�m�d�so�}a�C�ub;�;���dMb3���y�z�ۼ��uWU4y5=>F/ġ"���Չ-RW!�՗"$p\�>���S�w҄����vd������	4T���\�nƨP�ʱ:��ԝ�XLVt����G��5�&��p���P�#�|�B�X�g�i0\��.�gIt�!�����o����x�ҡ-�ّ�^ $� 'fa�#�i~0!�r�qU���Qv�EoO�؁'/B{�;4fx��V$�w�}MX�]y�y�3�˝��28Zlۨ�\�"ߗt$��6�iy��7I��XG��]�w9"x�g�Hz���MN����!I/�������A��1��+�W�Ń�I��-Nd+�A�+F�[���I\�wJ�G�����|�q<�_��s�֙���ƕ�*A�d�fWF0�M�J��@�WF;���.�P �0u��s$y���9����
�g�쎌�&���a�;�$y<޼e]]�q,�$X�刢0�]��	��M ?ؤ:�{��?�d���&�Q�.<�xN�[�����d(����I�ͭ[E~�ӵ(r7�l}�aB�g���B�
�I���^��*��O�t�!��6jV4�B��ٴ�� C�Q�+^�v�M�]�c۴l�&�j/vV_^{�^IN�f�w>{e�y{�הr�p�o27��e���im��1B"�A�`�=�ȭ^0E���^��0�$�ð��Tv��	�ʹ����?h���,��
��x(�i��/R�������	սL��$��ƹ���c�Xg�Yn��[_�����*�H`�~������w �I��!2,�4�+�-d��o�����x'=��O��(����<����+��!���8h��]$o8�(R�2�Ŋ�NE���5����A�>�xR�(V�RDFR7��U�z	��3�o�f���(�|�$��rÏ	�k�g�[�uQw�=+�����F�IQC`�%�l%zy�!jg�~m�Z��t�=Grh���?Zkܼ����Q�?������foȅ��k��4��s�S�,ii���5[��̔����'�u�X��@�v��~%BC�'y���xťwJ�G�����|�q<�_��s�֙`w7jH/g�3�G��+6Qk`e\����^�m�.4���2m�4�B��ٴm��ɅL�J)��e�O�{�h�� C���ŀK2���ƕo�����h4c�P�F~YEp1��t;��>��"���������X��1k��-��?O��xT�Z��5 
i�p]���#����k������CyC)ݼ�?E�~�#sv�RS�6���U��-|�v�LRu���$-��cLS��@�X+[%H����Ä�G�W8.+���W�dv��oTN!�������dҔ���Z��(��b=�i嬀֍�K�E�ө���x����8\l#�c�ۦ ���uN�;*�_��{M�бe���AP��=��;�n�dO�c����32��ӆo��*P�l$n�J[i���;��&͞d��M��V\�d	� 	qc�j�)Q��j8HQ��e�z�����,�W�B3���B[=cX�}��}v�_�j&��Ϻ�#Y��2�R�	��q'���y���4�CB��g��ۺ�D�͵SMI� y�r?�R�v~-}K�A�>�2�@w�?��?h��C���U�3�J~��k���k�[ݝ�B�W����k��)�-M
)#G�&���� d�":��p�T����pz��Ї��}I����#Q*b�6Ob���h+v҉����p�]ءVd|��()�T�~�k,9�? ��m�y���*>��$��� W�h�y��,-u��ƹ��t�d��`��'�BZ�-�a�Y�h�ݝ�B�W�ܴ����e.L*�d�,1X{���fz�}w�_c���\�+\�.��=YE��u��m�}�W-�W���E?��"�j��$�Lb�I�;�����k��\��@�u]�MP�T�%Σ��ĝ+����3J���|���s�44ȵ�B�B*��wj˻Z�zWz\ٿ�6�PG&XU��ѐaYR�B�\����K:C��<U_��s�֙f����h��y{�הr�R_ǌ� N��r*0��� F*,ƌN�jK�I�q������/f.������Ut�\��D��_:�!S�x�J�<�0|k4�Ż�&ǥ��a���F߸��S�Ȍ{ɝV�z����WN�d7!qzo_<�b"E��_'V��	��yO8S��%��3��J�:��n�&�E�aYR�B�\����K­[W�\M�_��s�֙]V�#9%���WN�d7!S�x�J�<�0|k4�@[�_zβr�v�������Q�^�� Fڱ���EC;�s�w{\�S�Ĕ�ZӞ�'�|,kW�F�����4�G�D�6(!rһpl�;�w����*H��M��FF�T	����$73���'���)Q��)���1
g�t�z�?�y)���t�%��	#�I�U�@B��rBWy03H��[.7|L����\c�;�^HUB����yt���w� �w(�
5��qD�KZ�����[�ƭM�R6�C1�f˾��S�d������m�I�_�k�8�ם��ɚ���ʈ�����)Hߋ,D���@�wR�� ������t^���\�}g��?`-ʂRcL�h�����WN�d79���'�!�'/2�%ͭ�=㜝�����E̒KV��	��y��Q�f<������E���YD�	��P�S�bN��E��锏��Z�� '����X,"�-��*1�#�;�����4�;��|B0F��#,k|2�Ω��!N�'�y�G