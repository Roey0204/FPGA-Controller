��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-@���rahZ����*��/}{�_@1������{S�������<�w$ɨ�h���G�m6
�DR���8�+I�S��n�D�N�����N�8t�>�Hc;��|B|X����}��_��t�ս߸�Z�C	�a1ﲀZ���dJh2-jwG�CUG@�t�k�k'v��ǔ{�q�%O���t����t�D�~w����+�#���]�0��mS��m%B����Ӻ��,Q�Q�?uG�Qy�����Q�Y�Bݣٳ���� [��(�� %����
�?<�곦���q1��B�ceH��.���s6�kk�`��y��&������i��0+�M��L,��.K��C���@J{�"F�6r/	�Y�B!zZ��۸9ߤ�Ha���3����!�L���!�`�(i3!�`�(i3���ue���!�`�(i3!�`�(i3F^I�i<}�sȸ�"rR!�`�(i3�4&8��z�[�X��ņ�3\SrXtN����f�%;.�J}��Ut���c�&��j�b�,t,�y�WW�W�ck��=~Ì��O�K�"��)�1������1������R���l%�odYǭ�%�Z[K�1��������;I6l��7�GQ�C����5�sȸ�"rR�· ���4���w0�DT��b֤�]�G�6���7��$�7��$EԔ	�8��6?���W+X�~{˕vC�|�ˏ8[$0�I�'�z��9���
�n|s�)>��!��<�ڒ�]X/��~�5:��fĝke�!�`�(i3J��+GP��fhH�{V�RDFR7�?D��׊�'�t+��u��^�ץ�7z��	.�V�~�-���\�>�/E�CԵ�_�*���d��4D���t���װh����t�D�R�WZ��@O���t��A�Pf�d�:o+'�E}u1�R�Ȫ~���		�X.]���}�W��� ���G���p�@OM.Ir��"���tc��=�����?�o�JH�S�Zt�(���b?(���&�!+5���Y�҃ڹ�^��2���96v_ �7�����T�٥��T)'��:�Jl
��Pn�߶h��Myf%���G�v���Y�p+�~��]a�{��>LTd��e�R��b�7S�����i�F��2�+g�@7��cؖ�r�M�?��	4�����wƃ(%��<'����Z"}�p����>�UKW�*�	S&&�s m�Ht���11
����}C9�S�+o���oBg�Caz�~�?���Bꮷ����A?�>�Q�k^�Á�)�o��.&l��ʩ�R'���=�\�W�EC�)�6-��~h�ӦI%}���/�çEF�)�]ܤ�1�G�Qc}y�����߫��Ѷm��Ǹ�vJ]�3�<
d�>��W����`�r����Fz�NK8�y �����<7u!�`�(i3f�s�J!�`�(i3NK8�y ��K�"��)�ul֗��|�!�`�(i3!�`�(i31������!�`�(i3&��潹!�`�(i3m�7�TG���^:��lFE�߇ç�b� ��Jײ?����!�`�(i3�m��7E��!�`�(i3!�`�(i3?������ޝq�~�[_.H P긭so3#���^�_!��� ���r�>��f1~�?��Ӑ����~�f h,��3h!�`�(i3!�`�(i3�· ���4!�`�(i3��J���FB���Շd��@Ő��t勪�i�/��{�P:tg��ݖ˘�&��Lӳ��{%_��6�z�
^��t&�"��+E�Tw�· ���4!�`�(i3h,��3h!�`�(i3!�`�(i3�· ���4m6
�DR�П�� j�L*կ`��%�����-���,���x��
R���eU<�������|[���HHi���~����Us��9�ۗ�蠒pP��!�`�(i3!�`�(i31������!�`�(i3&��潹!�`�(i3�����,I��Y7h�dČ���4�B��ٴ��s±���w	Qrk)F9�>�^W+X�~{��2�N��T$q��mKx"E&��� ���yoZ�P/Y�l��aLR����|���\X�TQ���EW�)U���a���C��iF�9�����$���y�VJ!���(�a��ܡ\{S�@g�(4������j��Z&��Ûf��O�.��+Y�B�&�%u�<��6u�G	O�V�g���ޔ��(p�]�u��.tƲ����%���a�>��$d�I�v���v,���h���ur�}w�*W+X�~{�ւ���z�X,mvvԩ|PM��!����E:v��M��n���/刲�Z��Utu⯃�ic" le�j�@���p��}K��f<�,=K�F~�?|�[_X��ˆk�=c�!8�Ԏi��p�7��Z鎬������~/[�� &He�ߏ=W�֯�^��N�&��?�2�1p�Qk�� h��ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08�tw:g�/�6=m�	n� ^�d�#2��0�DQ�L���EuZoO�=����'�ނ�ebÆ���p��'��aC�h�>�4����CX36-Q��ܹ��E!����梡���h�3��3%��׍����}0�st&���\�vūx`��:�֡�\�<7�X�e���V!���IÙ=�H�l��3d�`.�/'�����W;5B5Y+� �i7�sp>��=D3�OO�@I�I�z%��;5B5Y+�T�����N��=D3�OO~G��;ؔ�V@��n����&��J�f����t�Xx�s]���uC#����
p��#�IÙ=�H�&8���l�mq���)�:��j8HQ��e�z���V�RDFR7������`��I�t?�_��B�e�D�*�Y�p�Yч���Ҟ�+�����yq�_��x�s]���uC#���ج��iL�z��XP������<����Dg��y��tq�-[�v:v��I���w�����
�?<v�a�;H.;�i�����v@U?�_��B�e�D�*�Y�p�Yч���Ҟ�+�����yq�_���[�!U��#:a�0$2RX+�/�o�IÙ=�H�&8���l�mq���)�:��j8HQ��e�z���V�RDFR7��ᚌ��J��:sS89�*uT?�Х |�8�}7E��O��O
+@~`��)�j�����x�d��[04ͳ���U���O�8c�
p��#�IÙ=�H�&8���l�mq���)�:��j8HQ��e�z��͹sC�MP���!Z�M�I����&A��`�����i�t�<�<俇d(�D-rB}VGڝ�
�<��^�:�)_;5B5Y+� �i7�sp>��>9UW?8����V���Zy�>�@�מ�u��Ϣ�͹sC�MP7�B�J���1��b�,�MGuvh:a���(�[rÕ�)X�J�$�R�n"tXۓښ-x�]�V��o���\Sc��b�F�b  �H�,3�V���CS��*~�nzL͊�q�� Ky��:~d�_C�VJ����̕��W���x��%	#���H�	�q�@S%�����1&&��=ql��.�C$����}��yoZ�P/$zoRؗEI�$�R�n,�	�X�ɐk��@U8�JHn��z���G7�� �R���({&3�-��_�s*)F����Z�>)����hθ�|��{�r�\	��rR�Ɉf�=K����X���`�\Jg��à)��}�OV1
�Jzm���&��J����s��ވ�'��Ǵ�X�)Х��㵾�Fzjݭ�F���p� o��]���z��>x��F�\Mf���9��Y�{'%s��$z��"OW�fL�����20�3p,��ud�M�L�IÙ=�H�o��Je�����7!W�F��F�zL͊�q��b��~�U ��"�K�b��Ub�ۙD�^ֻ����XP���(B+r)��#P���P����ӑ7�\�<�(p�M�=�U� ���_�0)��ьu��D^�<�C!6�%��4&ݞ9��h�xm��.�3���l��q{�f��a�:&�>��s��f+c�.W¡����O�8HL�}mAb�+��XP���x^C�4�Z�U�C��z����1��t��YGQe�.-6�Qkw�<����SVcݧG �ŴP��Cn���}/�x�]�V���HN���McV��-H0
U�C��z���`�t�yU_� 4P/�W��[�&�pR<�K�q{�f��a�:&�>��s���7<]
Gxx�rDc�5��ja~��j.o�c�\.U1+]�!�;$��|��XP���x^C�4�Z�U�C��z��0�<��_MÕ�)X�J"��Q����%�8j�<1�9���9M�BϗHuLV��-H0
U�C��z��-p�Jj}Ѯ�/ښ[TJHn��z��G
�syP�.��:��z C��AͰ2��-��7�S�_�����c
�xG�M��ʚj�jY��Ig`i�ҋX����0�a1i~J����)cL�Z1~�g]�I���B��$ዶyHgb
�17��|B,����rY
��jP�9�D3���`4�E%v�~������]�!�����#e���5��(_]�Jg����-c �ЄW:zPCv����č�Y���S�)37J*u�v3���?_��PN��n�3���T�٥��T�xI{�X5�ҷ�������|���Aɘ%�ָkd�vu�Z��F����{l�f|�ό���.�>�j�gG�u����ov�~������]�!���#ʲL����M@3%�w����$ĄҋX����@�ڗe'�Lq���Bl$P�ĝ���1��P�߭�ҋX����@�ڗe'T���M0��s��]b_3#ڸZ鎬����v�Sq��}d���'��bw����$ĄҋX���� 
���u+�zN�����Ig`i�ҋX����{��}��^��}��~�Q��eHmgl���~O�Y5̹���>�Cb��{l�f|��rs�i��]g��u�x�s]�����*�T:�Ȯ��ߊ���&�t�),N�r=�}�{����0#��=��T��$Ю���ͤ	j�ס2��N�B~�Ǎ����+��|��].��'���Xw���,=3B�ݔ�]<�	����'rW��oV�dBmy;;���0��0��}���s��5Ǣ�{l�f|����%Hl܄�6K�u���"����o"x�ȥ��J���4�^U���	&}w|���!W_"z� �Q�c�C;=B>����}�v�B<��z��}�0z�cULv8�VWo�1�RR�,�*Ǚ62��˷���T�\ ���@��LĻu��w1j��a]��R���̠ӷ�&����>����Y�cӴ�"�6j���'��mr<�ҋX����0�a1i~JK>��{�T��p;��$�F#I�%�[���69[̰�&��YcH���V�^�h5��ٜ7t�}S��{l�f|�-�`��8�4n`�}�g���;�WC1wv�I�(��9�x���w����5I�E��p�)�3���i�A�K����
�?<J�!�Ӑ�JR����TD��ό���.�<��D�V��\�W�EC�X$�{�b�@IE�U��@�ڗe'	W��^$k�i�kL�5N�6�vg;Je'���Xw|�(���8��������)��[6���9�dMbZ鎬�����%�M��>�h$G�����=����(�
t��Y�{'%s=ͱu��̦�"�K�b��Ub�ۙD^�V]��}R�wX��y�J�#z����ͩ^��8k>6s����]�!��	Ǹ�y85�������&H�[&-n�g��U-�eJ�K� 3�d�����ca����{�/��6�vg;Je'���Xw�j�7���ᵉ3������|�z���o��W�j��6$>q��tm�Կ��TD���rs�i�����b���;���_�#:�N��u��_Ma�~�Ǔ8���/�L;� pf��i�!�� .�\q�K*'��(�
t�������2�b]�iz�f�؇��*�]��V-[q�P ڨ��S���Q�V�ɶ�w����������x[��H��z���8�ϑ��[���h=�������aD�orǟD�uiL${?���7γҬ�,;r�mR-AF�^ֻ����XP���1���*%��$�b��ev�~������{�OF8o/���Q]�.�Аs��J�.��ۦ� ~�p�tr��8`S�*���X���^ m�Z鎬�������(����5�	��]tr��8`S�*���X:�*��ܟ}mAb�+��XP��ș�\� ���Ӻ��L����~�pq{�f��a�sW��NZ�uw�@.�/wc1�
���D/:>mj	�Qiҗ�.̀�\�>�g1��< ��{��#�1d�v�~������]�!�����#e���d&���ݏ1��𠛕!��L��Q"��K,R��7��W`�����Z�Zn<˨	`�B)�}u��42�k����=g�?^<��z��}�צ:�)�<1(f}ظա�g��!ґ�E��w��RD�K 8�1�fT_UX�Y%/6��
����%E� ���1\U�_3#ڸZ鎬�����r44��ڑ�E��w���8<:XQiҗ�.�����k�f�[*$���6Ϝ�5W���s��s�!n}y���q���U�'ڐ�\{�ﳶ���y�B�M�5�Ta!;
=|s6|r[��bZ��b�Bv�~������]�!��%��rSe�u�heJ��Dv�~������]�!��	Ǹ�y85��r>?�W����/7R�%�T�\ ���p�N0��7Sx:��fl�}Yf�G�D(x���S'��%�u�p�f��$����_�}��Y!��TD�����%Hl�7Sx:��7�q��0D?e��{n)��G�D(x�듪�t%�a���̐�������� �������9�O���Òx8�!��N}�}���
8	*�?�*1�#�;�7��S�:I��w��,c�A�L'{Z�˗D�6���l ^�V]��}��kN8أ�>\��p}�	��D܂�A݁ؠː�� VU+I���]��w�sמC��_�2��+h���l`�M���-�uA^�Koْl��]�B9�θ�c}kÌ�s��X�e���V!���IÙ=�H�C�K2�n���������W;5B5Y+� �i7�sp>�%xI�ac�PƐt
׫�J��q{�f��a�:&�>��s���N-6�m~G��;ؔ]��ɲzL͊�q���������ӳ�Y�
�U�q��&�Z�>)������SVcW ��"vY0Jߺ�'n�^0o����SVcވ�'��Ǵ�X�)Х��㵾�Fzjݭ�F���p� o��]��r�p@iV�g,�5�Tz3�u,���W'���Xwd�n]N���ۆ7N1ƻ9��[�>�q�E#�UJ�#��Iam�D6�U6q��@%W�D�3����h������zL͊�q���� �Bb֊[
�}3���M:��2�7Sx:��fl�}Yf�G�D(x���S'��"�0ŏ�e����Ѣ�{l�f|����%Hl�dA���8��ea���||��/8'�L
�2�Ot�~�*�.iX�<�9{��!��{����t>=F�M���Yc)����]I�_3#ڸZ鎬�������i.ׯ�e>���K���6�z�
^7�q��0D?ߝj=N�$�<=�W�z��c�Z�H3=-��7�s|d_!�\�<��z��}�צ:�)7Sx:��7�q��0D?e��{n)��G�D(x��|�e�UTBfy���u\ع܄��� M�č�Y���S�)37J*u'H?�׳�#�,���Ξ7��G���C��g� ,f�?a˃��Q�0�	�A�����<��z��}�Q2�+�Yɗ�!����jT%q�#�<��z��}�0z�cULjaGkƊ~ݭ��%�x 7�v�ԯ�p C;8;���� ��[�����wo�A�I����dIϘ~Q��g&�<!�J�!�Ӑ�z��a7���6�vg;Je'���Xwe��(�R �p9F�d�<G� ���]��A�I���}��@�>��4���.����t���2E!^��@��1�@ �~)��*/�|�!���_- �v�j=U�h�]�vv���E�fZ@IE�U����S8��m�o�&i~G��;ؔa��-)�]��V+m�}.�Q�º�F����U�D�>i�ל�I�p\�WB��"?�N|I��`�orǟD�uiL${?�����>��yܛ�	��|��	(���zL͊�q���19TH���'�3�$ �#^�Vn�^ֻ����XP��Ȼ4�t=�j�.�/'�����W;5B5Y+� �i7�sp>��8"�@[�f;q�sɈf�=K�:���A0�	}�A�X5��_�G��Gq{�f��a��pP�o�0�CXL�\՚�P�S�bN֕L�����N��B�)Ybn���b���Y�I���^ֻ��)�cOKO&8_�0���@�p&ĩ+Ã��Q�0�	�A�����<��z��}�Q2�+�Yɗ�!����jT%q�#�<��z��}�0z�cULjaGkƊ~ݭ��%�x 7�v�ԯ�`�L�i���Jh���'�(���e����{l�f|��rs�i������*���ӳ�Y�
�Ɂ#�_���k�:�)� o]��8���/�^��/��L���WN�d7�בa��@IE�U��w�B[��lQ�$�k\_x���� � <�~��%���S��f�؇��*����
�?<1@�J�r�]��r/���梡���hV�W|�B�I:׷�F׫�J��q{�f��a�:&�>��s1�߽K}��[T�)���}0�st&���\�vūx`��:�� �����Y~��`�JKݗZ:���'n�^0o����y�]-X�G*.s�FÖ<^��4I^J<��R��"x��`]�n�p�'��-d�Ry��\�v�ȃ��X�\���e�Q8-�^\q{�f��a��N�J0���Uioέ���K�IE��;5B5Y+� �i7�sp>e�����1~��j.o�c�\.U1+]d�TpubMpIÙ=�HO 4v.Y��14�~�Xo��X�Ðﻋ-�����S8�E�qVf>&0I�=�H�&� LK�a�]G��wi�bZ��b�Bv�~������]�!��
ך��T�y��9/���`���6j��|E\0�*�W�ӝP�|��].��'���XwN�U�R��7W��!���{l�f|�ό���.�hM��{ �`o����;v�~������]�!��	Ǹ�y85���*�t�<�uծ/�,0=]^	�&������ *����h�(���e����{l�f|�ό���.ӂ����|�*3d��'�|��].��'���Xw�`��	��d^�qT�b㨵�֯��ҋX����@�ڗe'��.�f�8La���R�l�>D��(�
t�ژq���U����Q�S^��c-(���X$�{�b�@IE�U��@�ڗe'AKd��y c��"|�썥��9�dMbZ鎬�������(����l�`�n�>���/7R�%�T�\ �̈́��շ+���eq(1p <�r�\���ҿo�"aI��w��,)T{6T'8��������)��[68k>6s����]�!��	Ǹ�y85�Q��%s�@�zl���y���/7R�%�T�\ ��&M6^�Jm!�<��6�בa��@IE�U��z�г4>\��p}�	��D܂�A��W8ƭ�I�p\�WB����&�?�]�HB�ǇN��CY<Vf��?gْl��]�B�M:��2�$�R�ng~����2�|�]៽�q1�9���9M@�c�9�+x����"��Q����%�ދ����^ֻ����XP������'3�ț>�	�S�:�G~EiJ���ц��zL͊�q���19TH��>�ihbZ�������GJHn��z��r9�3��īO�8HL����K��zL͊�q����Ub�CP���{ƨد�p�L������嫃��Q�0�	�A�����<��z��}�Q2�+�Y�	q)�8
�L��W�eR���{l�f|�ό���.��6Ϝ�5W��Ig`i�ҋX����@�ڗe'������A���C�*�|��].��'���Xw�j�7���$�R�n�'��L�T�\ ��&M6^�Jm�{~�Ev�~������]�!��Zˎ�f+ոi��<�g�T<�t�S��{l�f|�ό���.ӂ����|�*3d��'�|��].��'���Xw�z%�ژ�(�WDv�b��h�Ӆ��x��h�6Q�7�0ʓY+��8k>6s����]�!���RQV�Ȭ�f�iC���R�l�>D��(�
t�ژq���U��C�k�j{�⳰��J28k>6s����]�!��Zˎ�f+� �߳G!�a�`��}��(�
t��Y�{'%s=ͱu���b�% ����ߪ��w������U2�~xao!f�	�Ĳb�M� �{��(�
t�ژq���U���i��Kqk�	(�´������TD���rs�i�V�W�+1M�`�"�X���!y(~,�a(􆿳�e�&���6�:���N3!�U\���<�����,�8��(�
t��Y�{'%s�h�v����}g��u"��*�ΊJ�O����	a(􆿳�e�&���6rJ�IaF�<��yѡa
��(�
t�ژq���U��޹ܮ�WB���k���8k>6s����]�!��荘�5V��ܤ�@�@yo�8�@I���M���J�ϑ��[���h=���D��F�omI�؝���B�]uo�s��X���n���Z[�ae!0�K�_3#ڸZ鎬�����۫s= O���t���x,pkXu��k ����ͫ��!n}y���q���U�s��Ę�5������:<��z��}�Q2�+�Y�y&��{)֍.�F�_3#ڸZ鎬�������(���n�Ak����
�u��٫7�v�ԯ�`�L�i�=as��9)NN�Y�N�rb<��z��}�Q2�+�Y� *����h��|���kJ�!n}y���q���U��C�k�j{����j�W���2uM�S�)37J*u��g���<c0�wg%c�_j��r�.������TD��ό���.�����v�� f�Lu�m�WT�j
�I��w��,)T{6T'�:���N3!!�[Oj8�6�vg;Je'���Xw�j�7���`]�n�p��h���o�8���/��
6�I��"�:Y3Iz�SŞ�Ӣ�8k>6s����]�!���۶$C�SC�(��EZ �:���Q���9�dMbZ鎬�������(����������TZ94��h���o�8���/��`��	����%n��WT�j
�I��w��,)T{6T'�:���N3!�U\���<�����,�8��(�
t��Y�{'%s�h�v����}g��u"��*�ΊJ�O����	a(􆿳����_k������U�p��
���)�"���R��� VU+I�"x�Q�jZ�|���!$�N�1z@�o	�Au�%]��g��xՉ�T�Ұ>D�c�lQKݗZ:���'n�^0o����y�]֡�\�<7�X�e���V!���IÙ=�H�]ƭ��&d&(C�#�7#^�Vn�^ֻ����XP���E)
i����$�b��ev�~������{�OF8��ڤ(������	��5�Y�w��~��Qg�.h���5�œ[�����p��/1Pr~�U�z	��U)���4�vZ�L��IzP���{ƨ���[AJ'&�_k�%w�_3#ڸZ鎬�����D�Kw���h`������č�Y���S�)37J*uc�A�L'��!�a��Wǖg3ȓ8���/��v.,-�{���[I��?ڔ��)KS�)37J*uc�A�L'��!�a��Wǖg3ȓ8���/�_�|fդ�n���i�+�WT�j
�I��w��,���|HH9M\��e���S���rB�6C�2��G�~�e�4�,���ۭ(��~T����z���Y��ݪF#.+����wU�ACctk��{l�f|�ό���.Ӫm��k�pN�By3��<Z鎬����r�1�	�0< �v�q�
�ҋX����@�ڗe'<��k����{l�f|�ό���.�@�L�q��(�
t�������2�8qTmI(xe�0
A���g�Lc!M�� �U1!ef����I���S��> �S 	���E�s��}�m�i��BԴ��ޅ=@��Ex!Ö�;�'���h'5S�)37J*u�t�H�U$�/D/}<�m*<��z��}�Q2�+�Yɨ��xvd�,�|��].��'���Xw�j�7��N��� ��V��_c�O"�Fn���H^Z鎬�������(���ȗM�+Ж�`�L�i�F̾0Z7H��6�vg;Je'���Xw�j�7��N��� ��V��_c��ڛ�R��'#�$�gZ鎬�������(���ȗM�+Ж�u��w[N7H9M\��e���S��> �S 	���E�s��}�m�i��BԴ���)d�ͥ�Y�P	dU�1Q��W��﹈�iq{�f��a�J)�!���[�j������z��� ܉���2Lg��`�+N��F.~O�,�=���P�r��ѝ� }o�!n}y��Y�{'%shM���VQ��W���:F�X?�g��U-�ei�u�r��F����U�<�]^�C��o�1t�"nF^�c�s�A��6U42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��Y7�u)S��r)�o�$C��c��(r���2r,~�oHZ��S�b=��%'�_��z�������ZI���~���U�z	��ߓ]�>k+;��5�k��y׽)N�[SV��˵��W�[4�	�}���^e@��V�i�I��Mֱ�H���� 5+� ��G�|��8��\n$̱̉���ߊ�,�'��.	&'Q����^�[��$*�¹�>D�� ��;����=IEw� e8�~�����0�H��OR�JO��V�RDFR7�h�Qf�����m���t���S�����ۄ؈��k�;4 e8�~���zR���bp;EK�6(��Mށtd؈��k�;4 e8�~���zR���b�W� D���>X[V��kC��8��h�Qf�����m��u&^3X���W��'LC��8����9&���"E&��� �����祎〕p�.��G�+-�q�,a��Z�q�,|�)�֢-du��~
�^^���X���v'�!��	�'�L��OR�JO����9x_�+���{�����w)�0�7��65�'�2%q{�f��a�eSܥOH�?�o>�q-7�� ��͌4s+�nyo�)��9��>x��F�\��Ɲ&���e�I\f"�	-7���J��ڮb�'���ߌ[R)Ms	[��c<+0.��Cҷ��eZ���hP*�g,�5�TzJV��šoLw8:Q�{4�5�Y�w���Q�`�B���B��!_O��Usj1n�1a�m�O��]�lEGV`2�s�f�6��5:xt�mdy�-��g���?�om��;���B3t�yL{�2{�=��E�Ծ�V���D/C�H��a�}8n�dY92"�f1�p,`V q��~�'�<�y8|�g�֐�o30�@Cq�,|�)�֑���w1�'f�wR�l�U�X��Ŏ.�/*��9J�]Sh�=�}�2����X+#��;ϫ�7�l�h�Iv01q�k\ ��e١g.�ե���.�U� ]��ɦ���2'\�d�����ca[�2&�;ϫ�7�l�h�I]����ljrk�� aD$O�x�Q�Q�?uG�Qy������(=2�u��s$y�刢0�]���,mxX=��uZ��הX{\�IV!"�:���l����R;5B5Y+�N�#�ɉ� e8�~��;�r"��[e�A`�M��V.�g�.�ا�v���}�{��<���#:B�Oy�~�R�&�����h�Qf�㷝�u!����7��=�B�z�\޳->��DV�RDFR7���X�A$(gKk��b�~)����n-Yg�yi��v�{�a�,.��/l8,�H����I��'��$�R�n����͛��W�c�'n�^0o��0I��I��'��$�R�n*d�c��n�b�a�JHn��z��`�B�92Y��^@!�PsgD@LM#��aPSp¦�5����`KW+X�~{�\���M�
`�t�啷�q{�f��a�I�4T�E��EMU�YG;] ,����a�� kF��4�	�}���^e@��VQi ��M�r��VYW\�z��j4��Rm�Ƈ��ݱk4# ��}��6���'n�^0o��3`r{�@~��6�% ���+a�G3�u]��;�LaP�'���ߌ[R)Ms	[����a�k���� v�D��qz�L<�������r���aM"��N�߄�4�X�)Х��Y[�P��)��\�v��N��V^���VB��z_��q�s-�#���[�"yd��N�}�g,�5�TzS�@/{�&ӧ�&��������s�����	)��59�M$#�fJ��<���6ɺN���ߙ߶h��M�k͝���:2�_]�5����`K�A���Q������;e5V�]C���[���?S�*���X:�*��ܟ���Gm_n��!$x�C˭oϨ�{�ś>���0�qU]�Z��L<�������r���aM"��N�߄�4�X�)Х��En:ъ�7k�%����x�ݠ�oY�1�O�vf���Wi����y�:�~%��;@6C�leKWa;.]�n{l5�z�}���XH���E>��V�Q4�:�^���A~��j.o�c�\.U1+]���H����XP���,#�N�MĐ�r�
���k�û&�l0�3p,����Ѓd��g,�5�TzS�@/{�& S�t����� �C��b���:� ߬����c��1���8}�Ͼ'���ߌ[R)Ms	[��l^V���
���*
�I��'�yۨ��~���CǍԽB�Z鎬�������(��＂��@ê�]���P�.�a(􆿳�tP"7��%�j)���������I��'��$�R�nL��C��&k-���h�����Hb�zL͊�q���es�1U)���\+N��&�L4⭦�����.��r�3�������r���aM"�������4�fN.�����?ׄ/�L	ACDCx��-��߂��g�K�
��$�~ȣ���XP���i�7��BQ���b�ǳ�LU�C��z��-p�Jj}Ѯ��.�x��W+X�~{�F(�E��p��+ᕮ��֫��XAьb2up,1�-�Y�}�ƈ�L�i����uZWC�O@�����K�Q����
�?<J�!�Ӑ�O���?�]�!���1����mB�8r\V��P?��������]�ٻ�q���U�pzl��a�V�RDFR7��/
����X?�WGc"�Ee�6;�ﻋ-���C�M��N�����ıψ6P�p�HZ5X�vZ��B��=Y��_�n������K�Q����
�?<2�,)�<xE;KC\�d�٣��c�A�L'M�Kc�I؆h��l7^*(��oD���g��U-�e�۴WLFo����|ՄT�٥��T�A��ˮ���nrm؊(��~����p�d~c�s�����_���&Y��V�c�	��}��/刲�ZT�p�n�ͩ���Z��]�!��	Ǹ�y85�L��0�͂=��«hj��I��Ba(􆿳�P��AK��hx��W̗���%��Aс�^�r2&����Z��beNY��;�W f�Lu�m�?�&͜�ﻋ-�����S8�r�:-�����`y���pzl��a�V�RDFR7����� �C!���'���Xw�����C����3��G�H�p0����ފ�:4*����X
V"i��rM���_��T���։�s/����R�AZ鎬����Ĺ#{��a'�<� \OYiucG�dd�����ca&��ࠅ�d�٣���,�JL���+ޡ)Ծ�͠�?N������
�?<���z�e��=Y��_<ͧ�:|�*�za�Hj���愝��C�3~	���>�Cb�d�٣���,�JL���+ޡ)Ծ�͠�?N������
�?<���s�6��N@u�p�VU��Jm�QA�Q* ��K�Q
�[�m�n�E�����Z鎬�������(���X�����llc�O��"X��[����fbK7͍��|��W&":і���#��%j�����x���s�KT�����bp�Mv�x��ﻋ-���`H�������Oд�( �#&�r�H�P�SyH���~}���+\�g��Z�&�Za
h�Q��<m��_���ݢ��d�٣��!�F8��_+H�]��>�YR��j5��C)���߾�'w��Mf���9��Y�{'%s2�ew��$�R�n��|��KB���`y����q����y}��c��v��P�:ݓ��E�� �߳G!"��zNt�NSx�lޞ��rs�i��=29��ab�% ����ߪ��w<��)�A�'�x9�5�L��W<Ʉ�n��Wlx�CzK��i�� La���Mw G,��LSx�lޞ�ό���.���K�Q	W��^$k�5t��v�Q3U�eT(�q���U�Мf�� �G�/刲�Z���c�}N�3%�}��!�������9/���`ދ2M�7���&��⬞g����[� hZ଻|�d�٣���,�JL���կ(����a�9���{��a]��R�Bq��jq:����@�3���3"�����r�&�O��p��Xę����'���Xwd�n]N�n�Ak���������Ll.�v.���ƶ�~b�!j��/��2���Qs�������>u~rۤG�#r,�-�_���c�@�l�ﻋ-���|P�������?xA4��Hݞ������;�9 �&x`rA���]�$z����fI�j�?x��������+w�7�Bmy;;���0��0��}�rJ�IaF�<J��d�X��]�!��	Ǹ�y85�����F�>Г������¡bfB��Q[�N|���OP�˟]��v�+w�7�Bmy;;���0��0��}�f ;+/��7I-G�]�!��^M���T�5xM����Qiҗ�.�˰m��T/��#���h����K�Q�B �n�6ӌ�Iۏ?�WGc0���x���"�Ee�6;7s�9���o�2�77�Eu��t�&6ӌ�Iۏ#���V? �#���	�KO�V3t;"i��rM�3���3"�ņ�a�t���EF�w*,Ht�b��<�d�٣��Y0����k�Dj��+ů�O��el���&����}l��r*�0v�y��| �҃�N�iP+��e�*u'���Q�@��߿@
9�"/����+�,M�}�^<o}?�0z�cUL���� @c�8���/�����w\�4��ղ�^��;,��*��� �`K�	����������n�&ʧ��Q���U�\���G��+��둵X�(Z鎬�������/�" �=�x�y��5m�xR_��GR�ٙ�=�T؅9;_�o�ȵ~pzl��a��yu>�� �U1!e�1�)��'���Xwwd�t�"��*蓱Wxi��U}t;#62O�a�P\�h�^��5�e`��9n3R7��)��-��g�SSx�lޞ����%Hl܀_+H�]��*ؐӘ��6�O�yc�������i����2ދ���A� ڈ�)�`b�\&A(`#d�A �W�rs�i��=29��a�����r���aM"��PǨ�o*� 7�v�ԯ�z�C���8���Lպ�t� ή[*%��JP�E��Y����|��Ay�'���Xwd�n]N�z_��q�s-�#���[�3��z�/��^�V]��}R�wX����K�Q����
�?<ТKH�{?����Y�Y�{'%s2�ew�ݧG �Ŵ
"4F��l���D��q&]W9	�׿*R�wX����K�Q	W��^$k�r�#;��B,J�j�FE�ﻋ-�����S8���{>�Ja�
��gl�4��H�������4�W�
�I�F��ޑ�L=�#�so��\�۟�-?�d���&����{ԕ�/�����jt���@
�ѝ<��6���P$��j�f��>0M�<k�lw�i}4���0�H^�wz�`h�?�15���{v��_G.B���uOܟB8�A��jeN�V�����٥����E�+'P2ӡ��,����|#^�Vn�B��מ�\P�O����X�e���E�+�$)�*C�8���EBy��J�z�3FN޻iai&���2nv���m���O�%� z����K�9y^6gV��Vv;�Oe�d�#�
�{�-������jb01
�;��S��y9Ez��}��H֞��� �z��w�����4L"炡t�8j�t�Y�Ij9���"]�ɋ|5��N���5�r/1ހĮ�J�z�30��G�$,Ek���J�j��v�x��W"����UK�B�%��ό�;�LȫԷ�/^�\MGl�<���{��ZT��6|�� =��_�Z�G�a}Cfx��V$�wpxR���B��Q"}Hi���#2�}����[��Y-��J��׍���o�B��^�H��7TB�7a	�����Y�
��3��X1�'�3�$ �#^�Vn���.,&	M��0�d�Sd��_�a���n�|W��ʞ-Ǆ36-Q��ܹ�q�i��@8���p�lő�4�`�+��t�Y�Ij9���"]�ɋ|5���F��S�%����&�M�s�F�:��8�^�.eO��q��S;gK�^~�U�'��gk=��[BfP3�e���b��M��Wv�'/B{�;4fx��V$�w�}MX�]y�Z��h��`�����o���c���w�L�R����*("ԛF�=���*� ��XLVt����G��5�On"WW��z&��y@���v���f��-/�J�¬��b����Lc�TH������7��ZΪm�T˚�Jz�0���je�Vmf��}S���u�����!S��cj^�+���Ã8�4��Q>�����=�>�>�(;��KX��ik���/҄UG�*"-M�O��~�/��J:f;[����˓#���Y!+����j�Ï��	p8,3s"-M�O��~�8(�#e��
LRi����o
��R/�[%씡����n?�q�Vٓ��(�����ꛓ�]�H@9�ݓ����6<p�W�4t8��?�Է�
��y��߾�'w���5����x(�i��/Rh�x#�L_�(D{ͬ�y�4������Q>�^2�����Vc2�����Vc2�����Vc�C0�M����B�|��1�@ �~)"���i01�(ZH4~��2�����Vc2�����Vc2�����Vc�����;��	�,G��q( �����k��S��S�h��|e|p�`&�厏�c�d~c�s���ݰ˄�ش@���&��~1E��}V��qO5�j�*Qtu�s�f�4\N��?	�n~�r%ӷ��Ø=%�MH�oO�'PP�~&�̵�6P�p�HZ�$����_w���O+k$�,P���ooF�!ݒ�롙��8��wJ��t�DY��b8!�ì�	jAKd��y c��f�\%�}���x$�;�6��Ѫh����
�?<�yǯϷm���\��E��U���}h��R�Q��=f׿�������!N�2��_:��y$[|�h���X �$�R�n�ĕ�dq�؀(�2�x@�����t��y�|�q���~�"����7Xa0~���;A���p�����|AW��ʗ&���MԲ���L��S-�����$þh���X �����R]Y�3�#�����T<�t�S�~�ch�B�_�+�)���&���/�"h#�)���w%e�3�!`�mLN��CY<½�T��+��������cx��=UW�l�l���XU(�a����ؽf���~�ch�B�_�+�)(�_ �¢~T� �}"���
wh���X ����
�?<J�!�Ӑ�f0{��
��y+M[K�}6��A�S�>�e�z���-k��f�	�����*�+Z��u��в}��B	�l������GVk�T�D�Q�(��s��8{�u�l��8��>ŔBU��o��ljrk��\O%�����։�s/�|*;q�rؼRo�~L$�������]�ۻ� �^�p�/�Caa��%3���o30�@Cq�,|�)��h��C�� �F���ꄓ��b&гm4���V���'�]ꅯ�j��\z��l��8��OT��)Ø����
�?<�9�x*�u����vj��'�]���-3FWҖ���	\O%������A��@���S�A}�k��&D��>�O��]��\&^�b'�û&�l0�3p,��~?%!���Z��0/zﴚ��I\CZ]��:f��;�46P�p�HZ�/?�?6�hF�Μ��EMU�YG;] ,����}��\>k�����W0TZ��7���">�3��x'�[�� <7S�*���X�#Gw6�E��0Tm5�q��4ȇc9 r�e�zf��7~g�[�!U���5��&<��iD�H	�����
�?<�09%?�3�1tm�/Y6P�p�HZ�/?�?6ר�`'֊�D0r➜~yٹ!5�j�B=?��FCC3Se�� ���� �C��|$T��!���o�8��14�~�Xo.ݰB�un����̧�f`�g�W���A`�M�7_]�4"m��򛘇n�Ux8
X	:J��Jt�k��T��kޏ�6j�"Hs���ػ!�&���\mИ|��,���לo�	�k��&D��� "̧�Y��kGQ��l�4��H���0�0�h��#g�k��cI��S}H`h2#25g�Ts��$���B�_�+�)(�_ �¢�R	d�jY��^@!�PsgD@LM#��7���lW+X�~{
h�q}lx"���%7B��0/zﴚ�T�p�n�ͩc�o�F=$����
�?<2�,)�<خw
�qNzx�s]�����!�C4@c���ė�P�"D0r➜~yٹ!5�j�B��}�m��V��	��y��f��h2�@�H�h��Z�2	[�d��x+a�G3�u]˴�����x�tƚ�e$+a�G3�u]+�u�G�k)�*C�8؉b�'��(�~��e�.5�����O��1O؜���z�h���D�3����h�>�0����ռ�ԡ�IQ����3�
+,I�20a���a�N�1�� ��2�����Vc2�����Vc2�����VcREBR�hHr��j�b�v��t��g;˥�b��a[q*�H2�����Vc2�����Vc2�����Vc2�����Vcɵ����6�pH�����qP��� ~��@���Wj��+��%S��P��}+801�)S��#)�& ܵz�"�st�^�O[H5�N�˼�v��j����&��J�eQ	�5v"���'sמC��_�2��+h���l`�M����Lx-�~x������������g�R�"Ì�s��X�e����]��m̽7a	����"���P1�߽K}��[T�)���V��ÑR K�R����Uܛ�	����$�c�=	d&(C�#�7#^�Vn��@�P��.�/'��"���P��ާv2ep.�����?>�Ab�_
�V��nyk��Q@�����8�4��_�G��G�����V1�=D�[ \��ݪ��fI�8f�Kuk;e�q��m�"V�40޼��r�p@iV�g,�5�TzS�@/{�&Zd�Zd�~��j.o�c�\.U1+]2��F�fsxx�rDc�5��ja~��j.o�c�\.U1+]���K7v�14�~�Xo��X�Ü3�^�XKS�*���X�#Gw6��>�u���g,�5�TzS�@/{�&qóf�ǡ-�#���[�"yd��N�}�g,�5�TzS�@/{�&^�V]��}�1�M]�6�k�#��.���t�:�6[��j;v��0�3p,�k�������(f���5C~��}����|AW�[5:n������h4c�=���� }hU��xz��osq�3�!`�mL�b�-G����� 5#�3��c�Ļ������rR��l����FZ�±��mJ^k��ô��Njr�Ú��k�VX��h�t(�ƺX���ϓ�S	T�	��p�q�����e8���Hmh���X �8�4��Q>�����#�FӃ(���e��~ж� ��%����
�?<�[gP�!�i��?Z4ZB,�D^Mp��$����_�!	b0�C}b�md��?�WGc"�Ee�6;���NǄ�{�#�	�����1p�Z�us�2���c`�V�s�]Ҋ��$�R�n��|��KB�4۞
�������U�p�6j�"Hs�g��Q��:nܑr�;V�E�S:]�c5���H����tV�������-�<�|AO'��ee=�4�_p��/v���5���Z@���L�U���;�A+b��}(���6�?�d���&��I&�^��7X�y�8Q�7��ʵ�<���(��h=��������(��x�l��15�r*Iީ�X��-�`V-u9�`�T�}��K��b�!cIh�{V/I�H/�v�6���l �-��f�&�L4⭦���;M^>+.���OϵA͆3�QH�ͩ/fP��_�����������*-�RԚf��Rm�Ƈ�hʨ}s��Zd�Zd�~��j.o�ѱ}����S�Jm gnt�S�*���X:�*��ܟDY~��;e5V�]C���[���?S�*���X:�*��ܟ�*��T�����}D��tr��8`S�*���X:�*��ܟ�9�4��'���ߌ[R)Ms	[��P�~�c��c��1���8}�Ͼ'���ߌ[R)Ms	[����Y`�^�kGQ��l�4��H���jȈ����Ӻ��L����:�k�;1?�[F�sp֟kh����aA�h�Ӆ��x��_���wg�W���'h�]^9����]I�r�B�,{�6P�p�HZG"{�e
Y�;���GU���|k��v·��\�RӲ�I�j�?x��n���Ϩ����t���s��Ę�}��U���)���w^J�b�=�P�K��J<W�f�ӊ[�k�T�"2o��3��	�3ַheJ��De��ڡ7oo-�Qd�|)3����ՀW�l�l���)���!���c�Ļ�+�m�r�d �~�ch�������l#QF�ky��.�"����
�?<�U
��ڌ�蜍6���e�|���6<p�W���^��G6���l �g��U-�e�-�L�=_8�c����sL]~ц>���K
�2<���9�m�w��v ��,�a.��!�s��P�����5������cjAڎ%�?��{P���B8���9����q�G��|�q<����a�����$�R�n�a��X�ktr[�h�_��s�֙�6�G�r-�k����-�����OD��vP��9{������Dʧ[
#���A�(QX?�>�����m�[0b%��e�旞f��T�"2o��%�������!�@�N�����p��R����K��aR�h���X �֯�ξ��k�<[*z����N-6�mmV�(� �D�R��_��֯�ξ�����p^�������
TF̾0Z7H��_�����
�od�6h�C�ˏ8[$0�}!v��C���[!����h���od���od�6h�C�ˏ8[$0��Hn����k�,������,�ǰ�AK�y�C�k�����d7Ud�8ձ8�#B%�_K:,�}ύ��c_C���-�L����)�u����D�{��/N�c�{�)&��{��!�T�.�w�$�^�QX��Rdo��W�ن��<�J�9��p)�i/j���p^���� o��u_��]�B�� f�Lu�m=y��lmb�?:��������8oOE&�O�Ep�z���}Ю�0��e0�?�����9䈔U4�$��;�\�'do�8qTmI(x;��|B8�}��F��O����4�)�Y�5}+�Z'� �Y�����
�?<��Ǽ:J'2�s |� *�9C���i&��R��x�s]���uC#����=z���j
?�d���&�D�;E��V���\U�����1g��d�����ca�e�9�2�����È�i�̠P�X:��"����0h�5e��8�ߧ\����W �-g	�X��d��S�!g�d���z��R�PP�_@Ų�։�s/�����"4�b~*��s�ݼ��P�v\�^�h5��A�$����@/��r �����%�������È�'�ߏſ�ټ�mˊ��ռ+���8�wFCR�7��։�s/�.�8�q�O;R*E���&�Ut�\���|��Y��^�h5���݄���'٥��gV�x(�i��/RŻ�&ǥ��a���F߸��S�Ȍ>`Β�C�3~	���ćh��g#ݼ��P�v\�^�h5��D����\�V��	��y K�~'&����p^����o�}�Xt��:J0e4x���O�?�轢2Ž;�F6��UQ@�������)�u����D�{��$�R�n�a��X�D�JM2�_��s�֙���^K��d\F��.��4x��}RBJ2�d1Z� f�Lu�m"���%v|(6j�"Hs�MR���I�J��X^��?u����j�_$�zՃO�߈Qm���ˏ8[$0���I�1(,.z3��o3���cli��7H�I�XHl�4��H��D-H�'\���|�q<��WV�#a��mJd��f�Ě��"��/f.��L�C���ea�Xi���y�����t���MI�wǺ�8Y)M���Fe-M�O��~�Ѩ�f?�R��֯�ξ���%L�#�R*E���&�Ut�\���|��Y�d\F��.��o(͔�%8n��뾦��X�H��Qߤ�N����
�?<�2��t6��N�g�c�`��rM�	 f�Lu�m5z�.TZݟ=�NM���ɛ�?ө�5ߧE4��rw�&�z<a��N� φ��<�6��̳#��d\F��.��4x��}RB]�QÀ��[5t��v��{����Ps_*�GqW�w��fD����
�?<~�l�>3��� |�=�b��<|)U�l��O�?�Ӌb,���T5�)�m"!�0�%�����3��/v���5����{�0����q�G��|�q<��WV�#a��n=�Z�@B��ї�ˏ8[$0�v'VQ�1_�p)�i/j轢2Ž;SQ$QW�b0���J�1��#���5l�qy�{���V+0f׿�������!N�m��n��&�7a	��������W5�\tCՌV�����,����_,�qo�,ܛ�	��������'�3�$ �#^�Vn���v_�"c�PƐt
׫�J��!��l��[�?2^�9,����_�X��-�`V-u9�`��	�����ɖ�V�̪ͭ,@�&>��@��H��pbn���b���Y�I��״��D�,҆��2��q&_���k�:]���9,�*#3���.�*�B�:N=����M���(f����j�ơ9��&@�E���+$nCe!0�K�r����h�ᮛ�ڥ��!���α�%����/�( [�� f�Lu�m�7���ŕ�T8i_�d�+��r�B�,{�5t��v��M;�E�iv�W�O�-�_���mATǥ��| hZ଻|�~�chXscr�2u��A�{(�_��Q�$G?g?	��o�cP��ym7��ҝ���1g�������;ϥ�WN�d7�\]�47����?t�+)�Lq���Bl$P�ĝ���	�}�Xscr�2upJV�ă\���q����� }v���L�C���ea�Xi�ݱ��/҄UG�*"-M�O��~ӟ�V�7lN�g����[�-^T/����f;[���e��@�����#����b����E�fh1f\����*�E��M@3%��H��	W�n�����%���3��a�����x��LN��v ��Lj�eSg��?`-ʂ��-�X��WG �����Z�[�U�߾�'w���9�2�L���Sӈ^t�lHn.��e��-
�8Z�&�Za
�����ھ	rw�&�z<a��N� φ��<�6�f�b E���6j�"Hs�MR���I��z=��ۥ�d���{+N�=ߓ���ܱ��K �?��}[9Ӌb,���T5�)�m"���F�tJ��Q�\��o�e/b�~u� U�X�l��%��)&��{�O[H5�NQCs">*���Lj�eS�������'�^����@[�_zβr��Û����ˏ8[$0�]�ν	��e�/a�=0���x����e�(�;#N�1�� ��2�����Vc2�����Vc2�����Vcv�iL�D
?X!��RS��uڜ3=�kM4v/���s�lIl��w&� 2�����Vc2�����Vc2�����Vc2�����Vc�?:�9�Ys�~f!�NE-7#еmݧG �ŴP��CnM:_A��k��u���?�d���&���u��Ѷ[?4���R;�9�2�L�+���\�RӲ�I�j�?x��n���Ϩ��IQ��t�Y���q�b�-G���G����@[�_zβrrZ�0m�\���>���=4�a��o��>��ʙ���-�7^Ya�:��H�D���Lxx�rDcѴ��B�66�i��ϗ=DUY=��ͥQCs">*�J]�3�<
��?��9)�r��\�ݫ�!�x���C�/7���L>Q;�im��9�θ�c}k���3��pg,lY�����y^Ii�M��oP�8��e�*���|��t��\nq��4�ca�(f����j�ơ9��&@�E�Ws�!R��p߷Td��#���~$�q����!��ZB����=�+K�����r�B�,{�6P�p�HZG"{�e
YR6�.�3��P�e�|��ooF�!ݒ���|kW�S/f��e�WDv�b��h�Ӆ��x��-�"E�}�����ņ�a�t���EF�w*,����n�#8�5z���GljJ�����v·��\�RӲ�I�j�?x��n���Ϩ��`��X~��������?��ًօP0��p�Q�@��߿@
9�"/�@��Flp�oN޼r[�z�Z<��zUD�3����h{d � J{?�d���&�W�!�
��i�!�� .���AOXu��w1j�C;=B>���h��ś͙��V���u��w1j�C;=B>���h��śa0��#���,0e�b��V��	��y>�w�`VFZ�±��m���*�N`v��%X��&���Ϧ)��|���؀.ņ�a�t���EF�w*,�}­]�Lb��[�-�0���E�+a�G3�u]˴�����x_��s�֙�������Zֱ5��4]�{�"�����{ņ�a�t���EF�w*,�AMX��QmL�x�3FZ�±��m���*�N`v��W#�����~45��<�Q+"�#�g,�5�Tz�o b�ўw�� ա>x��F�\�=�5j�˛|��a���V��	��y>�w�`VFZ�±��m���*�N`vR�Q�h�t5Az]�M�!Όg&W�w��fD�B �n�9�ǿvb���y�fJ\�/�:�Ȍq[e�-�l+7#~Ϟ3-��U�C��z����7��j�5ǌ��FK�~TP֣��݁#g�k��� �Q�c�C;=B>���h��ś�s���HAu��w1j��I����ТKH�{? ;��0��gBQ�*�Ѕ���ى�);"��PÛH�G:�g�]�zj7i�j��YoX�`�c�V��ņ�a�t���p
��9�GQDYR���g�0�u\=�~ o8�1�R�*���M�,������3~I/��\]=��"�ԭH���MO�/WOF;�Z宨¶J1�j"�A��"�Bmy;;���0��0��}�>9���־�f�iE�q�<�
�dSe�� �"���N��MY�5����;�
*�/�w� ��v���/L�^N��P�vJ}������eł1=S�B4�9T���l�FWv7�t>2Ϝ�Mg.6�kfF�5.]���ݾ-/�uu��ڿ$�)�vx��C�`�Bmy;;���0��0��}�f ;+/��g�镀��������ņQ�@��߿���A�U�u�;�����K��[��f����4�;��|B`���m򦨝-,e	�76��8�m�D�R�l��
3[ⱸ�ND[	��e��Ż�����r���aM"���Ig�{	#UEv�	��,���'�>�g;��|BĎ�|ł��@���:�ox㲐�a�A��ٞ�jBR,�á�?U�m[�c��1��;b��1�)S��#)J���l������$�~�;��Qz�#g�k��sИ�c�2Xy�WwꕶI�j�?x����� ���ѕ��J��!k/�5鎈���&��������h FS���Q;�im���M:��2�,����|#^�Vn�����'MB�I:׷�Fy�XZ@po��*���3m��U}�	�2�G�Ml\P�O����X�e���&qL�+.�/'�����WX�*�܁�c�PƐt
M� W��c+��k����`B�2�]�;f{(	,��.�����@	Qh���X �ݧG �ŴP��Cneɓ5o�0�W�}�ke�Ts
���!"����}���z��>x��F�\.��02��~�J��l�ꐘq?U�C��z����Ջ�/Cp�14�~�Xo��0���l�2q;H�-ވ�'��Ǵϴ`�-2c��ҭ��'���ߌ[��83�$^u������~��j.o�c�\.U1+]
n*�a��	h����Q�'���ߌ[R)Ms	[���$š���L<�������r���aM"��N�߄�4�X�)Х��=�\2�lFbI.����G�kGQ��l�4��H���jȈ����Ӻ��L����:�kg�m>�`^����S,د�p�L��������#�1d�h���R����	�m5�՞�ٟ�h���X ����
�?<.���6��l{��=�$����_�/S����u��w1j�C;=B>�y��[�b6����}N�M���$�~y��|�^4/��?E�l�1�ԀU�܄��� M��@�7��|���kJ��K�}i�e]y]�g��awf��!��ZBu��w1j�C;=B>�)3����ՀW�l�l���)���!���c�Ļ�+�m�r�d T���2�rۤG�#r�X{�"|Ӎ��5����'�)n�J�0/zﴚƮ�l��)8g��?`-ʂ���K7ή��B �n�6ӌ�Iۏ� ��*��HK�~8�zk�m1�H���W�w��fD�Ǒ�\�J;&�w��9�0��0��}�#b�j3�F�����ܥ[ⱸ�ND[C;=B>��\�����[H٠�X��?U�m[�c��1��;b��1�)S��#)J���l������$�~��Ŵ#����#g�k���ͪ	V	�4KCw.���6ӌ�Iۏ�=]92Q���B�װEl��9�4�~�ۉ�w;��x�l��1i�t�U��D5l�_�G��G2ŝ,\�=U�C��z����1��t!U$Y���7γҬ�,;r�mR-AF״��D�,҇��{|���?�}�h���X �ݧG �ŴP��Cn^�\���ĉq�p�F><1���*-�RԚfވ�'��Ǵϴ`�-2c��ҭ��'���ߌ[��83�$^�<ĘX.�
R��Ǔž'���ߌ[R)Ms	[����80���Z%ӗSu��z��j4��Rm�Ƈ��ݱk4# �
)�������4�a@�B%���O-�#���[�"yd��N�}�g,�5�TzS�@/{�&�<�?�aޑ�74i⯶��r�p@iV�g,�5�TzS�@/{�&rM$q�̅�	5�8aw�1�RR�,�*Ǚ62嫫�Rm�Ƈ��ݱk4# ���M3�=F�8�&��A6�k�#��.���t�:�6[��j;v��0�3p,���#ip��(f���˶HyNL���&@�Ex����MԲ���d��#�֢W�p�
ͭ��]I�r�B�,{�6P�p�HZG"{�e
Y�W�p�
����އ��&�nP{�B �n�6ӌ�Iۏ?�WGc0���x���"�Ee�6;��|fa��^4/��?E�l�1�ԀU�܄��� Mi�@�ZZle!0�K�r����h�ᮛ�ڥk:j%]a6��w%e�}�����ņ�a�t��T�b^ �%K!�Gr<�*���do��W�p�
͚�� Y�b�4!m4�UVu��w1j�C;=B>�y��[�b6W�����E��t�6��B�O�
B��$��~a$�B�X�"��ܒ��A��JrۤG�#r,�-�_���c�@�l��(M���9�c����U��\JD�@���:�ox㲐�a���)���IdiVbL� ��kYIį�a�y{�הr.}e�'�KBmy;;���0��0��}�<��WX��Y���jތE�b�&�q��ax��Y�L��x:A4bI�s�U�q �~k�%��x{^4��*m�~�޷Ζ� �1�f����y�F��K8v��"�����{ņ�a�t��|��[}����2��EN5L�`!|�l<�K�����W0TZ�gBQ�*�Ѕ���ى�);"��PÛ˻Q�0+�k��PHIO[9T���l�FWv7��:��~���vU�D�}�� �1�f����y������/��p�!���Ct�w#��@Ż�&ǥ��a���F߸��S�Ȍ�f����P��B �n�6ӌ�Iۏ�xA�)�Xy���!G6��B �nʃ��#�a,n�cqgFn�Ak���������Ll.�v.���ƶ�~b�!j���.Լ�;��|B`���m�^�>pg��	�}t>"�A����1sf�E��Q��-"�5mN ~Ϟ3-��U�C��z����7��j�5����z	�,O�*�ͳY����o�r%�fE�D�h�u��S/>��ᓺ�A��ٞ�jBR,�á�?U�m[�c��1��;b��1�)S��#)J���l������$�~�;��Qz�#g�k��	q)�8
�L!V�^���ȎS��|V�ؔ?%b*� ��~�8N|��7�'�L���E f�Lu�m^7]fn�c՝_�\�Zr�D�c��Q�Ì�s��X�e����]��m̽7a	����"���P��.0b����BC?T�<o�nïi�� T[��m��U}�	�(��Q|3�r�^K������О.�����@���U@���:��F�|4>��\-X�G*.s�FÖ<^�Ҁ��t�S��D5l�_�G��G2ŝ,\�=U�C��z����1��t!U$Y���۟D�$0-����G���y^Ii�ވ�'��Ǵ�X�)Х��㵾�Fz�������p����c��1���8}�Ͼ'���ߌ[R)Ms	[����Y`�^ވ�'��Ǵϴ`�-2c��ҭ��'���ߌ[��83�$^u������~��j.o�c�\.U1+]
n*�a��	h����Q�'���ߌ[R)Ms	[���$š���L<�������r���aM"��N�߄�4�X�)Х��=�\2�lFbI.����G�����20�3p,��x��δ�OUioέ����vЧ���y��,Zk�!7y�x�}�0�.�,�Mr]��F������#6�_���wg�W���'h_����Y�5X�vZ��Bh���R�޶(xʶ���5�՞�ٟ�_����Y��$����_�/S����u��w1j�C;=B>�y��[�b6����}N�M���$K��߶���܄��� Mh���X �����R]Y6]��m��bZ��b�Be��ڡ7oA!�䀯�'Ƶ�s�(���e��R��l����FZ�±��m>˟N�0D-O_�x�@��}-���?d����*�$����_�!	b0�C}��`Zf�Q�@��߿���A�U������*3���}������
�?<�U
��ڌ�蜍6���R��l����FZ�±��m�q1�i,��E�̂�(}��О�(ʙ��锴�;��|B���_|@k!V�^���ȎS��|V�،ܜ��hl��ם4Qb���T$�0��0��}�#���,�+� �9D^������¿-�#���[��0c(��<>p����ct�q�p�U��S��WV�#a���)�!�B`�� �U1!e��`���φ`Ldk�u8�Į�N��DM����p+k���HQْl��]�B/��v
���%0z���<��$�b��e�?��CG�����r���aM"��h�{V/��d�-ɇ<~G��;ؔ�Z�	����EYB]�.�Аv�മ#F>ͭ��Փ;e5V�]C��ؽMBW°��P'Q^|v���Q�cel��oW���r�p@iV�g,�5�TzfIT~�٤J��Rm�Ƈ$�pQ�!�s̽�_��z��j4��Rm�Ƈ��ݱk4# �
)����(�%�8��A���Q�� A�����>x��F�\��R�>�v^�E�Ή��Q$�@�xx�rDc�5��ja~��j.o�c�\.U1+]B�u���ASv�#�TH�N��}	��~��j.o�c�\.U1+]�k[�LD1�z��j4ݧG �ŴP��Cn**�8����>x��F�\�����2a�����E���˓k��i|Stߛ�mBp�S���E�������t�:���2F5���GݔO#�Z/��v
������aA�h�Ӆ��x�^�J�_-����h�}q�w�r\nȑ5�՞�ٟ�h���X ����
�?<.���6����X��H3=-��7����@�}z죹`Zf�Q�@��߿���A�U�u�;�����K��[��f*3���}�������R]Yp���Vh?�����=g�}~��d8���Hmh���X �8�4��Q>��5Zbz�Z��<�){:T���2�rۤG�#r�\���(.��--�7�Bi��?Z4Z� �7���H3=-��7��B�>�9}�����ņ�a�t��S����k��l#QF�ky��.�"cI��S}HbNzt��'M��WN�d7T���2�rۤG�#rUx��í��� �U1!eg��!�F;��;�YJ�� 6j�"Hs&	U��r2Qb���T$�0��0��}�#���,�+fO�v	B���� �U1!eE+� �ҕ� �U1!e��{m���}Ю�0C�Si����[ .p��A!�䀯��6Ϝ�5W��8	�+�P�܄��� M5�%!���;�*[�d�u��w1j�C;=B>�"�%|9�1���s�����h��N��e��b�ޥ��z[�g��FZ�±��m�q1�i,��E�̂�(}�-"?Ȇ�s��J?��N�)W H��YrۤG�#r,�-�_���c�@�l���=��s/B$8G&��zj7i�j��YoX�`�c�V��ņ�a�t��|��[}�GR�_[d����������Cᣨ*��w5t�}�p���� ��M��7<���Hn
V~$� �Q�c��I����ТKH�{?�7��|�K�B �n�6ӌ�Iۏ� ��*��H�E�;��S�UӇ�!-����,R?����>̞f�2-��������)�w��G*6}�{H�3)-օP0��p���Z۳
0.�
rQa��Y]�����u��w1j��I����ТKH�{?�Us��'p�-a�D͢�����.�x(�i��/R�*�W�Ǹ!2�͞nOYרx���*rۤG�#r���#�g���#� �߅�9�?�n9T���l�FWv7����хmF�wLoA���oq���--��w���L��m@[�_zβrrZ�0m�\��k^��=7�� �U1!e���aO��T�"u���t���ގ	�� ݧG �ŴP��CnM:_A��k�:N�si#�P�J�*T?�d���&����3 �rJ�IaF�<��*�J<l]rJ�IaF�<
cрp��sp֟kh��/ E�~ (6�3�SF�48�4��Q>�s��Ę�k+�xj������R]Y'�^��E9�����"�:9��HrJ�IaF�<S�	��<��k��qs{a�򖒒�����QS�	��z���n���u��w1j�C;=B>�v�{����A:��/��3:�u�jKBmy;;���0��0��}��`��X~��c��/�Bmy;;���0��0��}�<��WX��Y֊x���rۤG�#r�X{�"|Ӎ��5���l�1C��(�u��w1j�C;=B>�y��[�b6����}N�M���$
-��[ȴ?�d���&�u��w1j�߇V��H����d��՛� �Q�c���9x��i�H�֣m.�ｗ��u��;e5V�]C��%��Ob�|~qy�8:�d��$�j#�{D�A��R�3\�|���!$�N�1E��Zi���(%�9>��!E)ė(b>(>�}�����������g�R�"Ì�s��X�e����]��m̽7a	����"���P1�߽K}��[T�)���V��ÑR K�R����Uܛ�	����$�c�=	d&(C�#�7#^�Vn��@�P��.�/'��"���P���8�4��_�G��G2ŝ,\�=U�C��z����1��t�x'߼�p���+�M-/����S,���[AJ'&�_k�%w�r����h�ᮛ�ڥ��!����.i��M�R��l����FZ�±��m>˟N�0D-z_��q�s-�#���[�3��z�/����"X��[֗Q"t�����Jh���'�r�A�>$�!򆹋�I��&�A�߹�L:�%wk
F��.�
��吃1��v·��\�RӲ�I�j�?x��$�*�фXrt�&�m��2���<�(�A�߹z/�=�I=�t�+37/��Q�Z?�?\$��M��ݺ|��W�����ώM:��2�n�ڤ���[U�&�n������¿-�#���[�3��z�/����C_�!/XW�������f�w`�Ӫg[���+>g�m>�`^���t��˳���f̫zjI!JN��=ީa)�!��ZB��,�Ӏ(��[��B�IxoҢbu�ߞ�(ɡ�>�(}%@��7�����3�!`�mL�b�-G����� 5#�3j��dǑ؆�!��ZBu��w1j�C;=B>�y��[�b6����}N�M���$�@=���u��*�J�Ϸ���W�迿��!f�iBX[�� ڈ�)�`b�\&A(`#JU~akA7����ȗ,p ��Z�!3Bmy;;���0��0��}�f ;+/��c�%���pu����zj7i�j��YoX�`�c�V��ņ�a�t��|��[}�GR�_[d����������Cᣨ*��w5t�}�p���� ��M��7<���Hn
V~$� �Q�c��I����ТKH�{?�7��|�K�B �n�6ӌ�Iۏ� ��*��H�E�;��S�UӇ�!-����,R?����>̞f�2-��������)�w��G*6}�{H�3)-օP0��p���Z۳
0.�
rQa��Y]�����u��w1j��I����ТKH�{?�Us��'p�-a�D͢�����.�x(�i��/R�*�W�Ǹ!2�͞nOY��)Q��rIIksC-$�|���!oN޼r[�z�Z<��zUD�3����hY���v`?�d���&�����Y䆹��I��&�A�߹�L:�%��a���e�|���!��M;�E�����)��Rm�Ƈ$�pQ�$��ďn��Rm�Ƈ��ݱk4# �
)�����c�==�O��&�'ѝ�g,�5�TzS�@/{�&�o�^���p����c��1���8}�Ͼ'���ߌ[R)Ms	[��c��0�,ш��锴�;��|B������CUJ������wވ��hZ���N����o��Ac`��K�5�ba��O��.چ�$�û&�l0�3p,��ùd���M���Z�������1z#�Ǿ �� ڈ�)�`b�\&A(`#��IX��t�A�߹�L:�%�^�w���6j�"Hs�"iJ����~���.�Z�h�:�s�-רx���*rۤG�#r���#�g���#� �߅�9�?�n9T���l�FWv7����хmF�wLoA���oq���--��w���L��m@[�_zβrrZ�0m�\�z�ӛłMjή[*%��JH���A��2�����Vc2�����Vc2�����Vc2�����Vc��T=|ߐ�BB_m�g��t#�{�����^a ���N�1�� ��2�����Vc2�����Vc2�����Vc.�
͹U�5�X�W.���X;��P���P���Pz����[CQ��\�={"��sNw�%�a? f�Lu�m�/
����X�Lf�1_v"���'���mN4Y0]�Y,BM�Q��Q;�im��9�θ�c}kÌ�s��X�e����]��m̽7a	����"���P1�߽K}��[T�)���V��ÑR K�R����Uܛ�	����$�c�=	d&(C�#�7#^�Vn��@�P��.�/'��"���P���N-6�m~G��;ؔ�Z�	���$�R�n�6Knr�N/����L�zl���yB�cm��n ����TZ94���#��r�b�% �����e��7iӂ���(����kGQ��l�4��H���jȈ����Ӻ��L�g��Ԫt�b��r�p@iV�g,�5�TzfIT~�٤J��Rm�Ƈ$�pQ�9��j�Bl�14�~�Xo��0���o�\���a�U�C��z����Ջ�/Cp�14�~�Xo��0������CP��	h����Q�'���ߌ[R)Ms	[�����>C�1�RR�,�*Ǚ62嫫�Rm�Ƈ��ݱk4# �
)����Sc��6���N�߄�4�X�)Х����'��K�tr��8`S�*���X:�*��ܟq�
��sV$Q#�&ՠJ�14�~�Xo��0������&O�[
�}3���_����Mr]��F��i���k�bZ��b�Be��ڡ7oA!�䀯�Xu��k ����ͫ�I 	B��ˢs��Ę�ap7�L�	��p�q�����e���d����}$<N��e�|���6<p�W���^��G6���l �g��U-�e�����ߞ�)�XGGh���X ����
�?<f ;+/���a�{��t�����|ᷴ�P�ժ�Vh���R�޶(xʶ���5�՞�ٟ�Y&#�=å�FTZG|3�h���R���6���<W�l�l���XU(�a�<��D�V��\�W�EC�mg	}��h�6Q�7�����
�?<��X̖�	W��^$k�i�kL�5N�?*Yfl�.��c-(��96�O�n *����h�B�>�9e�|�3J��Rs����3�o�ll#QF�ky��.�"�:���N3!!�[Oj8�˵k�^�p�*��B��j��3�oU2�~xao!f�	�Ĳb�M� �{n�UYڕfC�(��EZ 4b�zvѓ�w7y�j>��l?
�A��t��#2��S���^RSŞ�Ӣ�PRۤ�P6j�"HsL_�4�8��CV�_!��e �������׋4>&:��Op�oP���kX_��s�֙T˷i�:�����
�?<1@�J�r�T�y<�N��ѕ��J�� f�Lu�m�n�@��N�������ώM:��2�$�R�ng~����2�|�]៽�q�E�u���tj`�;�_�2��B�>KUNo�^�8��!����29a���Qɑn&I�	~G��;ؔs����n{�>�	�S�:�G~Ei�J��
�o�${U��w�X�|0��X�~*�R���~�,��m[U�&�n��7iӂ���(��ʈ̩c��@�﹈�in�M�*:o�߈�vJVt�l�褻�sv�Fr�a��(f����j�ơ9��&@�E���+$nCe!0�K�r����h�ᮛ�ڥ	q)�8
�L��W�eR�l����%:x�6Ϝ�5W�!��ZB����=*�bA�Ë1��?��9)t#(@�$8�m�QKӲ�g����[����L�:�uծ/̫���Uh1݋��9�j��{~�Eh���R��J]�3�<
��5����'�)n�J� *����h,e(}�r�B�,{�6P�p�HZG"{�e
Y�C�k�j{�C�-VB�T���h�}q��������*�J�Ϸ���W<y�׀%\ f�Lu�m��v·�'�E�Jg�ˏ8[$0��I�tm0��f�iC���R�l�>D�iF'�� f�Lu�m^8��=as��9)N�*N/�p��3�!`�mLN��CY<½�T��+������%1���y��� �߳G!�a�`��}��P��hU�0��/�0,^8��-�H[����>�h$G�����:v�-�Yߘ/�o!f�	�Ĳ�z��"���0Yp <�r�\�w�Xb<��8�����p�D����13�3��ů� h�",oMG~�}�	(������o��W�j��6$>q��LO�k	q)�8
�L巋@*L��q.�)�l�dQIkT�	��<'����͓c���巋@*L��q.�)�l�d���{Y5o9�fP` �9�%��e�p���x�u���_;����X;��P���P���Pz����[CQ��\�.6e��H�Nw�%�a? f�Lu�m�/
����X�Lf�1_v"���'���mN4Y0]�Y��Ɗ[
�}3���_����Mr]��F��i���k�bZ��b�Be��ڡ7oA!�䀯�Xu��k ����ͫ�I 	B��ˢs��Ę�ap7�L�	��p�q�����e���d����}$<N��e�|���6<p�W���^��G6���l �g��U-�e�����ߞ�)�XGGh���X ����
�?<f ;+/���a�{��t�����|ᷴ�P�ժ�Vh���R�޶(xʶ���5�՞�ٟ�Y&#�=å�FTZG|3�h���R���6���<W�l�l���XU(�a�<��D�V��\�W�EC�mg	}��h�6Q�7�����
�?<��X̖�	W��^$k�i�kL�5N�?*Yfl�.��c-(��96�O�n *����h�B�>�9e�|�3J��Rs����3�o�ll#QF�ky��.�"�:���N3!!�[Oj8�˵k�^�p�*��B��j��3�oU2�~xao!f�	�Ĳb�M� �{n�UYڕfC�(��EZ 4b�zvѓ�w7y�j>��l?
�A��t��#2��S���^RSŞ�Ӣ��M��nq�p>W< |�;�Ojz�Qr�{S�$�:���N3!�U\���<��}O�Kz�4�b]�iz�?�d���&�0���v`�2�����Vc�cRq>ht�:���8��nQ�(L	º��	�cP2�����Vc2�����Vcy�Q��v�j����t��*��=@r�alb������t��2�����Vc2�����Vc��� �f��+�Ơ���r�j���Fu)n2�����Vc2�����Vcl��w&� !�`�(i31v��O�!�`�(i3:��B�Jz{#�a�!�`�(i3(�帿l�Lf�8�6�6a�}�_�!�`�(i3!�`�(i3���lx!�`�(i3��g�Έ9��n�7�YD�~O�h}C�_�Z���G
x�6�b� ��Jײ?����!�`�(i3�m��7E��!�`�(i3!�`�(i3?������ޝq�~�[_.H P긭so3#���^�_!��� ���r�>��f1~�O�xM�:	�h ���#� �-BD=!�`�(i3!�`�(i3���~>!�`�(i3��;�N�K�Ǔ�\=�����Y~]��0,Ѫ�P����5�(���עeqyȝ�No���o30�@C3)J}u�A�QOY��]gU��[�n!�`�(i3�7��$!�`�(i3!�`�(i3gU��[�n4.�����a>*�K��(�3Hzn��(VW�Q3��i]�������e-y���	�+w�`Y���2$6�sI#��9|�k�k�����Z������f�y@�.�gU��[�n!�`�(i3��g�Έ!�`�(i3!�`�(i3���lx|�G71�.;UW�
�2�8��o؏&�厏�c)]'SzȻz�� ��9�q�R#�S��ǟ��a��j����ZȆ���0`��WT�5˅������`dΜ��z(��$��=��$�R�nl�;�w����f����Z�וzj7i�j��YoX��0e �L�mW[�Ƶ\���L.���	W��^$k�5t��vl�0Q"Ob�&�q��ax��Y�L��x:A4bI�s�U�q �~k�%��x{^4��*m�p��vS�w��wv�G_WIR�Q�a�P�7_j��r�.��8b���6��{<v�/���jbPh<r�n��[F��K8v�u�1��s f�Lu�mr���l�7O��4'��7�OT�,ݧG �Ŵ
"4F��l���D��q&�t�>N�o���wu6��N}�}���<r�n��[�$*T`�̫��q<r�n��[�����/�z�X
3kZ�	W��^$k�r�#;��B�¶J1�j^aE,K9C���� �w��wv�G_t>2Ϝ�Mg.6�kfF�5.]���ݾ-/�uu��ڿ$�)�vx��y�D�
�b܉����A��V�RDFR7��
rQa��q�_O��������T�2V�q�Y�;�
�	���p	W��^$k��A��+�AMm?���e�c��n�cqgFz_��q�s|�3�d(]�/{��l��8�[��؁b����^�;��|B-��;qj���z� ��vOÉ`�B��5b��������`dΜ��z(��$��=��$�R�nl�;�w����0�0�h��#g�k��<y�׀%\ f�Lu�m�P�7_j��r�.��8b�����b��d� f�Lu�m��h;�ab���c-(��pa=ja=X����,�ǰ�I �9��,9��ҝ ��÷6j��1q[#+�m%V#2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�>-[1�p��}K��f<�,=K�F~�?|�[_X��ˆk�=c�!8�Ԏi��p�7��Z鎬������~/[�� &He��~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�'f�ٵ�J��ڛR��⾿h���l��q�J�2��C�`Q�%6�P+f�؇��*-|d{�A��>���K
��c-(���1RϦ�{8;�mVi�2�I�W�G���J�Q�ce��wRc��A�,��f3��uV�RDFR7��B�M�5�ߜ�7K����1�/!�������Χء<\:��{�ϥ��yoZ�P/;�y������,�p���>��yܛ�	��|��	(���zL͊�q����N�:�Pn���������W;5B5Y+� �i7�sp>7.~Ƨ����?2^�9<o�nïi�JHn��z��r9�37γҬ�,;r�mR-AF�^ֻ����XP���U�E�&�][�f;q�sɈf�=K����X���`����
�Wk;e�q��m;5B5Y+�T�����NG�2��o�7S�*���X:�*��ܟ>�V{\D���X���`���Eb�$3~��j.o�����i�]�!��	Ǹ�y85�>T
BFa@#G
WW�r>1�C�G��$���
G�|�!<غ��[��A���t�:��F{iY;��'n�^0o��p�N����.j�,�3*	��<�����j�b?u |�V���r�^�y4fCx=�a�#�1d�v�~������]�!�����#e���d&���ݏ1��𠛕!��L��Q"��K,R��7��W`�����Z�Zn<˨	`�B)�}u��.���6k��&�8�ҋX����0�a1i~Jьb2up,B*�U��9�����X)�K�b:GH�,�Y��?�N
���H��c�Ļ������r�!n}y���q���U����� ��p9F�d�<G� ���]��A�I���P5�� �-�"A�nTE�����R]Y�~�����ҋX���� 
���u�,���Ξ7��G���C��g� ,f�?a�+�zN�����Ig`i�ҋX����@�ڗe'��ՁO�#d�č�Y���S�)37J*uc�A�L'��!�a�&H�[&-n�g��U-�e��EB�v�hx��W��ר�>gm�Z�]�.nd�*�ۮ���1����)2����x�EyF�8ơ�@IE�U���2�77�E�ﳶ���y�U�z	��|u&��*�R�M���Q�2��`�3?RJ�/�?Ûﳶ���y�B�M�5�Ta!;
=1��A IHQk!��p�1C��'�ck�V�=��TD���rs�i�:�pdG��8p.������Y6�y!%O�T�\ �͎��ү3���, #3����;H/pH�����qg@ۼ���Y�,|3�L~΄gO�3f��*����f���,�L��;H/pH�����qg@ۼ��.s��|� �H��z���8�ϑ��[��2t�������?�z7����b���1�߽K}��׍����}0�st&���\�vūx`��:�,�qo�,ܛ�	��|��	(���zL͊�q���19TH��@���U@���:��F���V!���IÙ=�H�i�͒/e���@	Q�č�Y���	�I]����u/��R��@.T��^ֻ����XP������������m@�p����
��s6��\�vūx`��:�78�����,@�&>�;5B5Y+�T�����NK�w�o�k;e�q��m;5B5Y+���٫������ߞ��l�9�θ�c}k+�zN�����Ig`i�ҋX����@�ڗe'��awf���Ig`i�ҋX������S8�/ #O�)��BT�^��a(􆿳�e�&���6�L:�%N�Y�N�rb<��z��}�0z�cUL�V�xo�����@	Q8KߤW5�sH3�3P��[�Fc�k��`y�����b����蜍6����WT�j
�I��w��,���|HH9M\��e2��p-!]Љ������|��vt�����֬��g��i�U>.O���XJ�t21EL�́_� l�ߎ���#3���.�*�B�:N=�"���P�R��dˠ<GT�<PGc���7��Ǘ��*u�G�+-�=��a��|�U�N�4b��x��H����%QEIm{w�S� H����r��. e8�~��`:6`/�m���D��SW��Ƀ �Ώ��8�� e8�~���6��Z0��O,f�'}�C�=���a�Y�1�o<Z�L5RR������z�6�D�{�;�C�a�Y�1�o<Z�L5L�L�ɏg�wP�9�hE�u;Q��5�&�Jҙ�� e8�~���G:#��8,X���.�bI	\���&�Jҙ�� e8�~����J����a�i����\��O'x��.���]E��p�B�ݔ�]<̘�?8X8�Ԑ���%铿j���߀W~�s���!ns)��E�$B�ݔ�]<�����TZP��cul�ig"�SH��|�c˗��M��LG�IÙ=�H����Ԓ��v�1A��4�	�}���^e@��V/���lc�P��cul��iO\
Ǖ/Ds_���k�:q{�f��a�I�4T�E��p.�����Eqfv���ig"�SH��|�c˗�P�	�.��=�k2B]p�'���ߌ[��83�$^0��/q�1�9�j���B�<Vo�eo�μ���|�>x��F�\�=�5j�˛a(􆿳���i9����14�~�Xom�q�����&�;R�FJ.C�$4�	  Է�/ڍI� ����e�Iu����`B�� {�>|wՓ8���/��n(���˧�0z�cULY�ï��Jig"�SH��|�c˗��h���o�8���/�O�&�����'_@a���b�-G��F�i�w@`�d�٣��c�A�L'M�Kc�I؆h��l7^*�Թ��:�~�G4PN��g��U-�e�۴WLFo����|ՄT�٥��T�A��ˮ���nrm؊(��~����p�d~c�s�����_���&Y��V�c�	��}��/刲�Z����j���3��47��2V�q�Y�Hf�e\��� j�}8���Lպ�t� �(xʶ������C������H'";�0z�cULY�ï��J�iO\
Ǖ/Ds_���k�:��"X��[�{Ro�č�Jx9vyw���9^� P���&����3{K�BQ�tl��U������!�s����B�ݔ�]<�/����h#���m���bǣ�}|�\�۟�-?�d���&����{ԕ�/�����jt���@
�ѝ<��6���P$��j�f��>0M�<k�lw�i}4���0�H^�wz�`h�?�15���{v��_G.B���uOܟB8�A��jeN�V�����٥����E�+'P2ӡ��,����|#^�Vn�B��מ�\P�O����X�e���E�+�$)�*C�8���EBy��J�z�3FN޻iai&���2nv���m���O�%� z����K�9y^6gV��Vv;�Oe�d�#�
�{�-������jb01
�;��S��y9Ez��}��H֞��� �z��w�����4L"炡t�8j�t�Y�Ij9���"]�ɋ|5��N���5�r/1ހĮ�J�z�30��G�$,Ek���J�j��v�x��W"����UK�B�%��ό�;�LȫԷ�/^�\MGl�<���{��ZT��6|�� =��_�Z�G�a}Cfx��V$�wpxR���B��Q"}Hi���#2�}����[��Y-��J��׍���o�B��^�H��7TB�7a	�����Y�
��3��X1�'�3�$ �#^�Vn���.,&	M��0�d�Sd��_�a���n�|W��ʞ-Ǆ36-Q��ܹ�q�i��@8���p�lő�4�`�+��t�Y�Ij9���"]�ɋ|5���F��S�%����&�M�s�F�:��8�^�.eO��q��S;gK�^~�U�'��gk=��[BfP3�e���b��M��Wv�'/B{�;4fx��V$�w�}MX�]y�Z��h��`�����o���c���w�L�R����*("ԛF�=���*� ��XLVt����G��5�On"WW��z&��y@���v���f��-/�J�¬��b����Lc�TH������7��ZΪm�T˚�Jz�0���je�Vmf��}S���u�����!S��cj^�"w�Ln����	��#�WT ������5���֡�&Y��V�߯���s�Q��o30�@Cd�$�jz[�@!Xp��ݰ˄�ش@���&��~1E��}V��qO5�j�*Qtu�s�f�4\N��?	�n~�r%ӷ��Ø=%�MH�oO�'PP�~&�̵�H��2����Wa-�>���]k�kIY��oBd?\$��M��ݺ|��W�����ώM:��2�n�ڤ���[U�&�n�W+X�~{&���&o,>�*�B�:N=��(���M��oP�8��e�*���|��t��\nq��4�ca�(f����j�ơ9��&@�E�Ws�!R��p߷Td��#���~$�q����!��ZB����=�+K������g�$�G"{�e
YR6�.�3��P��q�����I���|kW�S/f��e�WDv�b��h�Ӆ��x��-�"E�3�!`�mL�b�-G��i�w��[5l�q����T��Wjc��,��ѤN�#���������2�W�8�q��T"��9�m�w��[�!ܥ�)�û&�l0�3p,��~?%!���Z���}?�N�*�9�m�w��b�-G������b��V�RDFR7��3w"��R	47�2���Rm�Ƈ$�pQ�$��ďn��Rm�Ƈ��ݱk4# �
)�����8�B����&�'ѝ�g,�5�TzS�@/{�&��@��)��I�-�A`�MοQ+rZM�H@[�_zβrE��g�Hbk���3B <��g�^^�xS��~/���jbPh�[�!ܥ�)�û&�l0�3p,��ùd���M���Z���}?�N�*�9�m�w��b�-G������b��V�RDFR7��3w"��R	�h�����6j�"Hs�"iJ������c-(��=��n��MBc���i|Stߛ"�st�^��'l7Ӱ���i|Stߛ"�st�^�[��r �%aWp��.�替��+���<j�_D�E��Y���{b�#�Uioέ����go�+��On�AN�.p�"z>O�q���<�{�!���"����d�#(���L[��وH�{�G̔�1s���O�Y��#~G��;ؔ��Νd[�*Ac<�p{�^���\�}����
�?<=�+�	�;rYپ�#��}?�N�*�9�m�w��b�-G��������/����W+X�~{�A`�MΈ�BT�^��a(􆿳�h�Qf��?Cb4!ޒ.C�$4�	��^e@��V��Ȫ9ƹ6j�"Hs�n�Y f�Lu�m��M;�E:1�7!p�"w�Ln���*v����t��r^1B�ݔ�]<�H �^P4��c�.[K��ml�;�Zݛ�\>n�Mw�/ϙ�v9�����X��o��4�$
���"Dʱ���4���Ewj�,
O���|��dq�e$��C��iF�����޹���#1�(Vc�����D���y�	),�Q�^�� \����K�w���)��)�*C�8؉b�'��(�~��e�.5�����O��1O؜�(�@�~v�]9Zb�;�ģ�4!d�B�
+,I�20a���a�pϣ�و�پ�&�̶�i�y�q�L�P�G������ޣA�лmm�����"`cI��S}Hd/S4T�eGz 	~l<`,9�H�W� � �<;����`B캝>+�W�^���\�}����
�?<��5���-B^b`��q\��������ώM:��2�,����|#^�Vn�����'MB�I:׷�Fy�XZ@po��*���3m��U}�	�2�G�Ml\P�O����X�e���&qL�+.�/'�����WX�*�܁�c�PƐt
y�XZ@po�	s��NփZ���0�lf�'��w��y�j\+��8����Y�I�����k+ �6����?�y)��{�!�e��f�F"�:f��^e@��V�苢ѤZ��h;q Hd�ٹ!5�j�B�)�p*��W ������D�J��s�;�9D�Gۥ������F���9�@Zd��`�H�&���1DV�H��~ж� ��%lsσw�kz��ՁO�#dh���X ���){�ו�T8i_�d�+��r�B�,{�a���ʔv�sNރ���Â�&�V���do��Tǥ��| hZ଻|�~�ch{�#�	�����1p�ZߤE���	�����U�p�6j�"Hs�MR���I��u�L��������w����'���F�