��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���a?K���J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-���տ��ê�Y�o�:g �C��A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD��aC�h�>���SW͟��W��x[����Ȅ�\#+��S��3��3%��׍����}0�st&���\�vūx`��:�֡�\�<7�X�e���V!���IÙ=�H�l��3d�`.�/'�����W;5B5Y+� �i7�sp>�2jL�K�B���.D7�GV��F�-���o��C!T*�q���U����Е� �7Ê7�E�4'���Xw<b��&ɛx�����4�b�k��g���7fj�~���3PS���X��u��(�
t�������2�=�����R�S��q�P ڨ��S���Q�V�ɶ�w�Q�41�&��~�I+����R#e��ds�H��b�^5J_�>�q���U��ȓ�iӚ/��Ϥk�;��|B}ø��y�w���H1��@�	��hN�q;�ǔ10\p c
N1�V&�����O�qTkή�Ádo�dvAg~�rk܀�#��˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F�;�sB*�1v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	��]���������ї4�z��pU6�M�S��2�{��΂DЫ�5�E-%Jn��ɧ���7�)a���%}D������h�br���lpda���\��6m��B��${��?�J�Z��]�Kt�E*�#�,���ns)��E�$�v����ox3��vC��Z�G�a}Cy^6gV��Vv;�Oe�d�#���!��@HW7��ո\����8�L���9���D�K�X�Re�d���L$�ѸT���C6���$73���'���)w�i����0\p c
N1�V&�����O�qTkή�Ádo�dvAg~�r{m��<�te˩���.|��f�ͣŗ�:���+"�9���B�I:׷�F!���H�v�!���y �谝��X�e�F����To?��m\Ӓ�qܛ�	����%��1����ї4�z��pU6�M�S��2�{��΂DЫ�5�E-%Jn�p�+~� �yKYQs��[�|�F��˱4���[�jDG|��o"� ���I��Q�yt�G��Eׂ̎�WI�;�_�	�t쩖NUD60L�b�J��@��y���Y
���^�.;��L�O<^��`Y�F�����I��#��
Mc��������=��:p��C��8�@��y�.��3��pƼ�+2!n`�pάYc:�IX[��O2 7�,�)�C5�!f�f�2�c���w�LnXZh��\����L�Y&8���p�lŕ��W�������9��~j5��Fo�P2}�).;��L�O#t����n��]ߺ�`@ZWH]�+Φ���0+C�yk;� N��r*$7�门Q��Ȝx� uŤs���Pg�H��
E�j>Pݮ��?��yxP+�L��k"S�	�C����xQ�n
V~$�Y��Z%][��"��z�"�d�q9+t�}Ż�&ǥ������3�$�Y�2�&��*��MH=|#����ڂ�x(�i��/R���������V���S��3Ah	)ޟ!N�'�y�G