��/  J��S���J��S���J��S���J��S���J��S���J��S���J��S���J��S������ ���h�k��$�J��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-
Ү��p7ŉ�x-�)��\y���{�z�ox�!P���b6�')Ri��_�
h������a�;5B5Y+� �i7�sp>1�*_��h_�
h�'ʯv!	��;5B5Y+�T�����N1�*_��h_�
h�Su�X���;5B5Y+�0�T��:1�*_��h_�
h��!n�x*4�^ֻ����XP���3�Tt
�w�}of�O��p�k����\�U�q��&�'n�^0oO,�����5����`K:���K�n̙z7��(�Ԕ��~��'n�^0o���{����I��'�S����cܙ��u�X����W�,���Op�ե[CF���y7�5����`K:���K�no*��\MI2#H:�d�TpubMpIÙ=�H�{	�� =�R���c&;�/��V��WB��	K�U�&��9�Sca�&'�'n�^0o6��U�x���5����`K:���K�n̙z7��(+�}�Ҳxh�믳��"5� �S��Z ��d���%�a�A��CN�vs����L ��xQ7��y��Vu��s$y�4�Dg2^��I��'�S����c��2gF����Z8{�):;5B5Y+� �i7�sp>1�*_��hjOhi��ȫfc<�R{X���w��|��kVU_�E�I��'�7w����w��Z8{�):��W0i��^g��F����%�a�A��CN�`ѽ�N��}:�E)�F����@��zL͊�q��K��e�m��0nZo�j���
,H+�Ӂb�9�f��W0i��^�A�hA�@O1�*_��hjOhi��ap���
)��;�}�u��s$y�4�Dg2^��I��'�S����c��2gF�����ͧ���Tq{�f��a�P9b����%�a���錜c��=�
>��$0�"��	֧�ǌo�9񶺸��_���׿k[Ai����@0���u��s$y�@�~T�@��5����`K:���K�n�Z(J,��*|��:\��^ֻ����XP���3�Tt
�w�Ocm�r�?���0�i_@#�8u��s$y�6��ܡ�.�5����`K������*|��:\�+��CY�E2�e�.�
11�*_��h�����T��u�{��2.��p��3�̘*T	6�'n�^0o _xB�I��'�!f_\eN�g	M@�����W0i��^�A�hA�@O1�*_��hjOhi���Fϴ��hۃ�T���|��N�p9:O�I��'�S����c��2gF���^�iq��;5B5Y+�.��h��u>1�*_��hjOhi��U_�8��oْ�h�R��|�����j����I��'�7w����w®^�iq����W0i��^��7H��R?1�*_��h�����T��u�{��2.��p��f�\�=����\�v�ʁ�t+o���5����`K��m���L��Lv�
�Sx��=֧�ǌo�9񶺸��_���׿k[��㴀@=��EĞ��W0i��^��ѫU�1�*_��h�����T��u�{� u�WA�=��,�Ⱥ[�IÙ=�H&+��/����׿k[LTaL^P���}m$��|�����j����I��'�7w����w���T���s�"5� �S��f�H?͌4s+�ny�Gz�SQbʛʇ_�^�i���j�b2o�`Q�zL͊�q��e�[,E0nZo�j�:|'4�e�2��J�h{o��W0i��^�A�hA�@O1�*_��hjOhi��T����%w�|���_n��Op�ե[Qq
˟6͌4s+�ny�Gz�SQbʛʇ_�^�[v5(�#~F�Qm�JHn��z�����͉͌4s+�ny�Nh�`(��OX7|��,��s����Op�ե[c������͌4s+�ny�Nh�`�sS���j��,��s����Op�ե[Qq
˟6͌4s+�ny�Gz�SQbʛʇ_�^�i���j�b2������B��\�v�Q�����͌4s+�ny�Nh�`UN��`v�*�����.u��s$y�6��ܡ�.�5����`K������&��C�<A�������92��|���{�.��y͌4s+�ny�Gz�SQbʛʇ_�^�[v5(�|+��	�]y��\�v��1�bC/Oy͌4s+�ny�Nh�`(��OX7|�0���J�J�u��s$y�6��ܡ�.�5����`K�������L��Lv�������92��|��HRC["b���%�a�A��CN�`ѽ�N���� ���;5B5Y+�Ȩ�� "�DX@^w
��j��A6�]���`$��ؔ��/��:K�vV��7$��Q,�!<�/�P��=�﹈�i��W0i��^�A�hA�@O1�*_��h�����TKR�Hr/�@��١9�G~��ڹ 	�"5� �S�"� /`�j��%�a�A��CN�Tk�.�E<��Cm��'�M�il|*_u��s$y�@�~T�@��5����`K:���K�nbAUL���K�"E+F�ؒ��UeVP�?��{	��A��@1�
Ү��p7ŉ�x-�����[�/�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'���?���ʢS����E@��<��W��k�۸�y�uZoO�=��1��AN��!�\#Ƌ4ͭ�'p�@�,3_�f�_8\/HiO���L�~�$�d�?�%�7P��T���\�vūx`��:�VŤ3+���;ۂ��IÙ=�H��p�ӷ�Sw�����3ݢ�2HL�JHn��z���-&�@_�!�7@�7ы��$��9��}�.ޢo�%�D9U:`?cq=}��r�#�87��8���#2�f����[�/�-������|��%v&ͩ?�>�ɻz��wSx�lޞ��rs�i��|,�xh�G���);�y� I�Û�]�!��	Ǹ�y85��P���Ԙ��ł�!r�dN�<@Iv�,.9�������? �mV�
Z����q{�f��aƑ��t�ڣ��-)��_�|��vt��p�/W
�'��27���A��B�6l}���C�4��3n�Ĕ^ֻ����XP��ȽFBcl�����6~J�I�*ط�c�zgV���gVk��1`����lI�35m��\�v��+e�Z~F]k�4.���a�����-��z�/ �,Dp��u�����h��uR�p#5�tҗ�^��lI�35m��\�v�[�w�����=MZj0��iK��h��P�Vf 'R_���GFS҈�l���D�V[�>��{�|��	y��~�f�'n�^0o�h{4N'��	aQ�� xS4�q���-���^�}������jK�P�nH�]��i��� �;5B5Y+�T�����N���y��lD+h5�u���Ͻ�Zı\G�+��C�W�2$S��Ѡ�i�L����`4�E%v�~������]�!����͙IS��⿣:�d��{l�f|�ό���.�wZ K�Ϋ�v�~������]�!���&7χ����n����$�_3#ڸZ鎬����Ĺ#{�����݈>��}U����B*�2���u���d���� 	�� <�`�hE���Mz��;��ҋX����L$�����/�{��U��+�����E)S��,2�����^���@�d�_C�VJ����̕���(��h��+��<ȫ� `�r�d�=i"}�۞h�G��L/��!n}y��p�VU��J}\�=���(bY,?Z1~�g]�I���B��&���a�%�j@c�rn7Zմ#&<D���l[�!'lBv}��q��N��f�;�>)�'^-�G�0_3#ڸZ鎬����Ĺ#{����>d�pāea���||��/8'�G~+�3;��\���\��k�zph5)�� ��i���ӹ2��c=�_RBD{���p�9z�AR�v�~������]�!���\B��Vp�E-ޕG�g��$y�z��eU�e��������Dg��y��tqӴ����s������"|����N��� 	�� ��I�}j����CX�ҋX����L$�����/�{��U��+�I_�=0<��,2�����^���@�d�_C�VJ����̕���(��h��f�<�K6���x��B�����_��K����č�Y���S�)37J*u�"��ȝ��h��� ���ѡ�e�LZ\^ �@'�ZX��<����L�Y&j8x��l+��DL).��\1F�5�ͬ8�.��č�Y���S�)37J*uc�A�L'�f?S��##�'�\�ge��T�\ ����S��G9��f1�p!!v*!��u���d�Ӵ���)�jj���|}��3�G��T���93����R��Vj�'�B�>�9���9�dMbZ鎬�������(���kk�ȥ�S�}���G��Yʬ`�f��`y�����䫦.iK(�au|�I���B���
��u5YM)� �G��U�
�d�3��AR�:�Q�%Z��;"�,Y�i�#��Ig`i7G#+��Q2�+�Yɑklb\�PQ(J�i�5��^:��7+\򃘴�WT�j
�I��w��,�=4�w�ͳQVia�Y�����c��7��+H5(��?��6�vg;Je'���Xw���e�Kfx��V$�wo�1�:��L~΄gO�3f��*�����th��#*��1T~��3x���� �sVp�Ͱ����`�orǟD�uiL${?������{�c�t}ܹ�~*JHn��z��r9�3���.R��ª�E"�'n�^0o����SVcm�������RثNTu��s$y�����SVcl��2G(\�[B�����'���Xw���'���E��}� �l9��9?_��=Y��_�0z�cULL�֗ul?�T�\ �͘�f��p�b�z'hۉ)r�k��)�νY�T"�W�F��F�zL͊�q���^v��<f��S��E�j��
��c��1vэ��wL�\�HlZZ���!�Ѐڋ�?躷Eښ�ez�JHn��z�kČ���Y�� л���&_��q>��s#�9���&���.R�%�N�YE�WzL͊�q��j�|Su����geEq�l���j��k9���'�L�,Ot�������Y���h��崸{�|��	y��~�f�'n�^0o�C�~��j�4�aY��`ս�B���dV<4����;{ۤ�&�TF�jK�P�nH�]��i���{�|��	y��~�f�'n�^0o�h{4N'��	aQ�� xS4�q���-���^�}������jK�P�nH�]��i����{�c��ai	�z���XP��Ȇ· ���4���6~J�I�*ط�c���>s˘�ؓ�_��C}�K�
�4l��T�#%��B�ip��{l�f|�ό���.�$���H��č�Y���S�)37J*u)T{6T'��osq��|��].��'���Xw�V����t��k�|��|��].��'���Xw�����C�;R�<kQ~w���~��ݏ1��𠛕!��L��|��k<�<�`�hE���Mz��;��ҋX����L$�����/�{��U��+�����E)S��,2�����^���@�d�_C�VJ����̕���(��h��+��<ȫ� `�r��Y�Ȅ�f�;�>)�~�`�0��|��].��'���Xw�����C��Z_�� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j����H��[n��B��X���WΓ�BD{���p�պ����u�Q_�}{KS�)37J*u�,�JL�������d���J�l�]�Jg����-c �ЄW:l�mq���)�:;o�����G�̥}�ߘ����N�[վh��[�3c/��!?V#$~@!<��z��}�<ͧ�:|C���m9�/Ɨ@��ݏ1��𠛕!��L�ވ���ۭNJ?�s�C�,����&�2 �����&G|2-m�Y�Ȅ�f�;�>)��5�g��|��].��'���Xw�����C��*��z�)� ���ѡ�e�LZ\^�e���Eы�`�M7Э���j��S��^1���k(�2��c=�_R�*�b�m���K����č�Y���S�)37J*u)T{6T'.?-��o@�e6qR5L�/8'�L
�2�Ot����F�2�v����oe#<�ފ�R0�z6UDu\��-������K6jT%q�#�<��z��}�0z�cUL���gM�6�!�u��އ�e���3a(􆿳�e�&���6�;�x����~kE#z��eU�e��������Ӟj��s �׊�8²u�8���=ON��t*�[P{C�#^؆�PĔ�5������:�TD���rs�i��=29��a��>�\Ԍ�m��H�^��"X��[�`�L�i���(�M�D�bó=��!��L����犷��r��\Uo"S�!jw�bD�h/O����Ҡ��Nv����V�/�בa��@IE�U��@�ڗe'�klb\�PQ(J�i�5@F��a~��/(�wT�בa��@IE�U��@�ڗe'�/H `����,}��յ��lY��qq/8k>6s����]�!��荘�5V��ܤ�@�@y��a��l��0xCv���p�3	qA�ý�ɮ�a��t�?,���w�F��cK��{�tn�a�N���_�\�Zri�;qGܒ��(~D�2h���X �7�� sz��woT�c��v�l���Ҹ �gO;\t�j-׬�o��y<�ơ�Ǉg[����Ĳ����l��2G(\�h���X �o�u?Yɲ���woT�c��ƽ]dN�4�Z;��1Е�j��2K�q :u>m\f���<UI"���4�b�%Y�w��Ǉg[�����S��7���� �Ǉg[����)��;��@��[
�}3��*���1����1�pi�3h���X �{Ē�����B��+��р��U�cE�i���f{ �$��`[��8�Q��jja6JMԲ�������BNC1b��%���۞h�G��w�O�r�e�7�gI��<�`�hE�n7^��_�۞h�G��L/��7�gI��h"r��n7^��_�۞h�G��n�oS����ߗ�H���3c/��!����L���e'��ǩ��b�N~�+��Ecc�,�[`�7���c`e'��ǩ��>F�q�u�>��Ecc�,�[`���ׁ(B��
,�U&�o~�H�C[c����8�0��$˘-�������K6��%����_$W{���`��:BY����^�i�����m�q���z�n��9�n,]Q�yfT�9������h4c뻖*����u��z�	:�h���R���M%��3+�7�����L~΄gO�3f��*��������[�/�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�yߪm����Y�{'%ssA'���?���ʢS����E@��<��W��k�۸�y�uZoO�=��1��AN��!�\#Ƌ4ͭ�'p�@�k�U��ʧ�V���,\ަ�It�i$�$[���ɾ�;ۂ��IÙ=�Hb�����K2�:�5q{�f��a��4�6�tڬF
��[lD�����.(��"5� �S:Zot�{> ���{�c���
È!�Z鎬�������(������˚�9��9?_��=Y��_�0z�cULL�֗ul?�T�\ �͘�f��p�b�z'hۉ)r�k��)愥���ޤ7��;ۂ��IÙ=�H�42_�'
�7eUshl~�Kϯˏ�K�������ܭ�'��:�^��8�m�\�=�1p��'n�^0o!��0ך��$��o��}M��`�ܜFS҈�l���K���qb�%Y�w��;5B5Y+� �i7�sp> �d�n0�����9X�O� �VI�:iZ�Q,��\D�ш���g������E��Vib�%Y�w��;5B5Y+�T�����N �d�n0ϙ�K4`����j��I�:iZ�Q�K�3X"��6�!��w.�4iI��d����|	q.�q{�f��aƩr*�^�	�<�6�Q=S�W�$E5<4����;{?^�Z��μ�P,Uw��ZmM��j+���0%ђ ��zL͊�q��J4����(���H�Q���12\p�G�iAL��K�~����.j�,�3*)���U�7P��T�<��z��}�Q2�+�Y��\�6�(�_3#ڸZ鎬����N��q���$�7P��T�<��z��}�Q2�+�Y�>�~I� �_3#ڸZ鎬���������4nNt��k�|��|��].��'���Xw�����C�;R�<kQ~w���~��ݏ1��𠛕!��L��4_�;��	�[%�lM0�u�Q_�}{KS�)37J*u�,�JL�������d�?���Qz�]�Jg����-c �ЄW:l�mq���)�:;o�������{���_�G���;�Ζ"�љr1c�,�[`�9+��d@���{l�f|��:2QYeƈ �-u���k��H'�񽂳B*�2���u���d���=A�2�S|���f?��� <��U�-�R�so�	�C�d�=i"}�۞h�G��n�oS���|��].��'���Xw�����C��O��"�( ���ѡ�e�LZ\^�e���Eы�`�M7Э���j��ᶨ�8�U�}{����@��WΓ�e'��ǩ��b�N~�+_3#ڸZ鎬����Ĺ#{����Aدo�zea���||��/8'�G~+�3;��\���\��k�zph5)�� �T�5B���"�D<�4_�;��	�ya0���Uu�Q_�}{KS�)37J*u�,�JL�������de�0��`v�]�Jg����-c �ЄW:l�mq���)�:;o�����p�ǔ|�b������\�����	�-<����Z�E詄ҋX����@�ڗe'.?-��o@�e6qR5L�/8'�L
�2�Ot����F�2�v����oe#<�ފ�R0�z6UDu\��-R��C������Ig`i�ҋX������S8�����)�d=1Yih��Ïx�x�>J�g��U-�eP�����b#���w*͛����6~�I���B���
��u5YM)� �G�=O�@���<�S?�Ϳ[�3�~�2	[~U3�&^��0� �8k>6s����]�!��	Ǹ�y85�c�l��o|B���x}S8#K_���8���/��dQ֮��R8�Ņ�~L�e�LZ\^ �@'�ZX8�5}7�ɐ�����A�H��E<lKZϖ�L��6Zr�j��7P��T��TD��ό���.�6��GJf��誆�J��������/(�wT�בa��@IE�U��@�ڗe'X5M�����,}��յ�o��C������9�dMbZ鎬����+��4{��M��y��I�sVp�Ͱ���@m��0�&���#�{�0;�}�^��w
����W*�XөF�;v��8�v`A�2��cN=�vAg~�r��{� u�ll�Yɍ�ȩ��F}Z�J_m��nB�ft�3����dL�o{��~�,�lRo+&J�E<7�����|�"ya�= �'�Q��f/�����JDW�%-C��o;v������Uq���V�PQ����h=��;���yW�B��c�Ym̚�s�M:]�Idr�xR$TP�W��	]�	�"Gr�v�� 8��P�>	��� ����˂�i���o'��#{��pj;x7q�|��ł!��1�ϚPI?ȹܹ���8�v������=+XR/ v�DiT��Τ�<(���t/�)5�(���{�eV��0�dy��8ۦ� ~�p��71>ڨ�/p�ַ�sA�jLt��/�U&���#k� �SMӱ���즀e�E����}�cϮ�(z�/}=��_W7¤d�<�f�Ģ� ���y��U��?܅��Xm�>��tI��l�b��i:+���F��K9�_��(�ʵɿ�&Pp��.��Y��m�^��1�Ey�(�LV5��B�\��4����h���E�&����f��jv�!d*�[��
ņ�&�&���#VW�GaAO�� ���V����&��0,�]��s����w����:�y��9�\#���8ᅧI��v�u�%"��a/�S7�<h�����)`;�+7��u�+�y�ߝuL���I��p���	[⍒��Us������,�2�(������b�_G�KҨL*�ї�>EtГ��lW
맻�_g���U�QH7]�����_kzO$8�� ��b��c� e8�~��(-��xsF�o��ǵ�ڊ�X3U�J,���b�,�����e�V�L@��$���uȚk�&���hڦ�	m���N���[��=�<��^~�y���uȚk��f���[�q�_�7�vw������A���f[`�-�z��Fk0�Y�{'%s43u�R��va�Mf��.7�\�x��}���G��t�B�Q$d��^3�I!^�V]��}��ł�!r��V�e^笾8�4)r�=��{Bhv�̙z7��(�C��E����'n�^0o:WB~�z�nF̔���>�\Ԍ�j�O���⎢r�
����X�$S �;)��ơ��SYƒc�������m��Z��h/����� ���c��_�&��9����H�~�u��8
��}���G�99�����ת<����9��r��]��5��f�4
�Ǽ
�����g'�Y�
p��#�IÙ=�Hn����2�4w��S�Cd4�\��� �F�S�:���3*���Ux���� ������/2C�6ⰺ�a�%]��g�ܐU��\�7խ�W0i��^��(�̠A�V���߃�'n�^0oޖW�/�
�^�=�Q��M:��2��h���_��{l�f|�ό���.ә�ՠt9N�σQ��Z鎬����=���ޒC>.��ކH�.7n^^'p�@IE�U��@�ڗe'!����b�&�b<X�'���Xw�j�7���˷���T�\ �������>�F����UR[Q91��ۆ�p<����I�p\�WB���b<�B뿒x�=��[,OV*�؂9� 4
���;*�,���^�=�Q���fɂۅ�M	���x���yyZ鎬�������(���R��F�D�g��U-�ee�@Rv����my$�N���Uە��`ZjS%;��k���'���Xw���ؑ�
@��,�m4S�)37J*u�,�JL���
����v}S����,�<��z��}�<ͧ�:|��ΥT�t�U��1<<ap��hٳp�VU��Jm�QA�Q* �R���&|~�i��ft��]�!��荘�5V��ܤ�@�@yȻ�o�?cq��c�7h�	}��A�"�V�RB^�&!��t��\#+��SЫr�T���>:&���W0i��^������:N�ŀ�9MpW~�b���{ �-ؼ�6@���c܉y���VD�m�F"� 4
���֧�ǌo�9Մ�:n
eoq�������*�9k��/����@IE�U��w�B[��lQ�$�k\_x���� ��٤#8,ܶ��ahC��PT�bEl���"��ْl��]�B�M:��2�nˌ�!5�_����
�z�8ے�os��zL͊�q��W��{z'x��ū��!Vi#@���%&E����T�Ӕ@t�iap��hٳY�{'%s2�ew�~�G4PN��g��U-�e��0v�p��<��Q�'���Xwk�~m�nM���f��k'���XwL���a�G�;ɾ��Z鎬�����R5�8g:ؓ)�L���Y'���Xw����#񯢝{l�f|�ό���.�L�6�k��ҋX����@�ڗe'ѡ�MI�#I��w��,���|HH9M\��e���S��JvW�����q�@���N��]�aՒ���D|-o�Z��beNY����X�	�l��f1����]�!���1����mͻ�0� �]`�Jt��ﻋ-�����S8�~3i0'x̙z7��(8gS��;��T�\ ����M��a�Oo���+��t��P� �M�q�Z���'�W8�7ՙ�V�-7��ﻋ-���C�M��N��dP�ɨ��1�Z��[B�����'���Xwa'�<� \nJ���	��٨�.B�ﻋ-���C�M��N������(��&*3�,u�Mf���9���q���U�pzl��a��y����Ig`iZ鎬����Y�V��#q���ɨ�ML�9࡯�d�٣�����6>���]�B��[S�7P��T��]�!���1����m���!�����Ig`iZ鎬����Y�V��#qt,�����Ig`iZ鎬����Y�V��#qb��Q�dt [B�����'���Xwa'�<� \c��`ʗ�Mf���9���q���U�pzl��a�ӫ�$�߇�Sx�lޞ�ό���.ӜM�q�Z����z��T�KH����
�]�!��	Ǹ�y85��~�g���` �f�N�g��U-�e5��e6²�\j�>:�,1~����[�Sx�lޞ�ό���.���K�Q��C���_����k�]�!���1����m�\j�>:�,Om�u˼Sx�lޞ�ό���.���K�Q:o�>W,���Ig`iZ鎬����Y�V��#q3Ψ���=��~�����ﻋ-���C�M��N��X�N���XTt���9�&��=Y��_Q2�+�Y�V������o~�H�C[Mf���9���q���U�pzl��a�E4��8���W�+���zZ鎬����Y�V��#q��9
c����'��]�!��	Ǹ�y85��_3�i�GT�#��+���������t�&��SN��6&� ��=Y��_Q2�+�Y��������3O�3�r��Sx�lޞ��rs�i�LZLø�ʞRW����Z��T�\ ���|.�Tӏ�b1�t��ts�vbp0�]�!���1����m��w����9=W�玞���K��pzl��a������	���嵓'��֔�����>^�2�����Vc2�����VcREBR�hHr�A��5�V�����w)К��g: k��2�����Vc2�����Vc�t����?Պ@9)�A`Ј*/��W�v����%��v��g�L��:�WT��8�|��&��x����b�G���l����ʎ��J:)�=f��F�fU���[W~L��?�Tm#����Xb�r�I �۞h�G���',�K/{J }dx>3-���t�q9캧xӍ.�����{�T�ؼ�n�B�'��D�Mp�=n�٠��f�;�>)��-oO$t�&k��@f�6��	=Q+�����3c/��!�����g*�s��I�G��L=���;�H���ou�QR)o��b����;�H���o��և�GI-��N���xf���2�����Vc2�����Vc�m7���ee��j�5�>�[L��2�����Vc2�����Vc�$M���l���ۢ�x0/�*�>��"�$-���`~[[z�'K�$|��]4�lWh0��p���Z��xGj/*V�z�{,�lѩ�{�F7�'�orǟD�uiM���	�fl�Dߠ˨�R+d�8Dѕ��e����������T���0�|U�.h�#nn?l×n
9�.��_��C��N�'�m���1�R�M�&H���١9�G�29a���Q\f���<Uȫfc<�RE�AE|��GݔO#�Z/��v
���p'��'ׇ(�x6�'�rc����8�0vN^!�a�]٣�2e�tV��	��y������3dF�N���O.�^����,�,�}v~�GO>��-G�r�6���`ѽ�N��}:�E)�F�t|���^���\�}�!�c6���V���Y')������Ȩ�,\ަ�It}�0�.�,l/u���!�'���UV��H M��� i�A�/8�M��)Hvl/u���!�P���sA�el$gS��:���K�ne�rE�*o.:���p�+~����f�[ۻƆeu��<̮Z;��1��be�|Y�l�r"�'���GݔO#�Z/��v
���p'��'ׇ(�x6�'�rc����8�0vN^!�a�]٣�2e�tV��	��y^J'I�.�o8'�ij�@��t�BLf-C�C=rGO>��-G�r�6���`ѽ�N��t������lH_���U�߈��<�u������RͩɮpƆ�H����4H�W������������z��,S��l�ǈ�J�_�Ǉg[����o�oߨ��o":�"eġpǆ��J�`�Ӽ\���L>�vHUHN�ʯ$�4UBQ�/�*���jš���:Q�l�H M��� ��
,H+���~�O����/��NO�l����m�=�er߮��h���_�!��ZB��e�s���񱽽&O�c����K"��rQ�4噃,Eۍ=��w�[l\� C4���IJ�.i��ܰY�̄��&|��}��m��6�,t�#g�k��lvЃ",3�@�'2��A6!p�-�ْl��]�B/��v
���+�K=�Jᬉ>:&�h���X �7w����w������<�l/u���!�P���sA�el$gS��:���K�ne�rE�*o.:���p�+~����f�[ۻƆeu��<̮Z;��1��he���O�(�$(�ʭ!7y�x�}�0�.�,y��w_8h�y�,������KA�E�#>�����U�p�6j�"HsJ�[z!p�ũ����˃�ud]�kݹ�I�4~��J�6���0rk޾�Z_�ʇ_�^�[v5(�ͭ�'�qj󸤀hZU�߀QG���ɮpƆ�H����4H�W������������z��,S��l�ǈ�J�_�Ǉg[���ȉ�k�־/R���kE��a���b��]���;��d;��f��2R!�u��އ,),U2�CM��G�j���&"���vIh�e�B>l�2��!f_\eN�_��Z�0����~�;����ɝ\�!2A`ZjS%;d,��s�J2����I;�H~w:��Ps_*�GqW�w��fDud]�kݹ��u+�r���s�Y.��A
�7�$G���s��DX@^w
��=��E&�����L?�d���&��kv��'DP��ju�Yz��J����ܣ٧�\�T�q�>�YŇ=�er߮���^��oF�v�മ#F� �gO;\�(����>̪���$��@�Pd	���~)�iI�
���1vs����L ��xQ7v!:Ӽ��t��ж�﹈�iǇg[����I�u��Zn�Yh$W�x/EI���āsp֟kh�ҳ�	�(�ω��t�}Qhh���X ���K�����(M���9����,�ǰ��>,����S"1�(L�w�X�.BO&�Ƃ۾�F!�9I�4~��J�6���0rk޾�Z_�ʇ_�^�[v5(�V��/N�^���\�}C�V�4�Xa�,h�V�|��-q�ٜɮpƆ�H����4H�W������������z��,S��l�ǈ�J�_�Ǉg[���ȉ�k�־/R�L�q�G�	
�̔�}9MpW~�b�B�GQ1{��S����c܊/��8muS���dWk[�W*e/
Y��g�'�鶴���;� �gO;\(��OX7|���( 	�Gb�GݔO#�Z/��v
���p'��'ׇ(�x6�'�rc����8�0vN^!�a�]٣�2e�tV��	��yX���)��2&�Eq�o�'��>�w&�����l�p����Ŭi�O��<RʉGO>��-G�r�6���`ѽ�N�����C�H_��s�֙��ճ V���;MC��q�����U�յk`����&ߓ�J�X,��x�l��1i�t�U	
�̔�}͑!/0�D��nj��L�C���U�":�"eġpǆ��J�`�Ӽ\���L>�vHUHN�ʯ$�4UBQ�/�*���jš���:Q�l�H M��� ������0�s?�2)�/EI���āsp֟kh�ҳ�	�(�ω��t�}Qhh���X ���K�����(M���9����,�ǰ��M�J6C��;MC��q�����U�յ��Xƥ�o��h���j�_o�'���ޠĀ�=����+'u��ɛ��`���u�{��C�*�����`=���[���Z����jS���L:-�z�Ry۾�F!�9�V���Y')������Ȩ�,\ަ�It}�0�.�,l/u���!�'���UV��H M��� ��pR���J�h{o0�|U�.h�#nn?l×n
9�.��_��C��N�'�m���1�R�M�&H���١9�G�29a���Q\f���<UU_�8��[` ������/��NO�l����m�=�er߮��h���_�!��ZB��e�s���񱽽&O�c�����d�.f~銐D�_g��h���_w��Yy���(1�G#?F:�}�7&����Ŭi�O��<RʉGO>��-G�r�6���`ѽ�N��)&%�����;2����Ls?�d���&�[k�'*�FRO�}�1c�K�7R�;@��{�E�x<��J����ܣ٧�\�T�q�>�YŇ=�er߮���^��oF�v�മ#F� �gO;\�sS���j��\�y:�_�]מG�u��t��?��CG��>�\Ԍ\$⨹�2H�Q�i���IK��m�F"&[�Z�{����m���L��Lv��0>� 9�/EI���āsp֟kh�ҳ�	�(�ω��t�}Qhh���X ���K�����(M���9����,�ǰ.�A���dΣ�J�o�C�%tJ\a~!_�YPj3����.-t�O���Ŭi�O��<RʉGO>��-G�r�6���`ѽ�N���-ޢMr���1D�牆���Z����jS���L�.-t�O���Ŭi�"ˎ��E#PA6!p�-�ْl��]�B/��v
���+�K=�Jᬉ>:&�h���X �7w����w�ޔ(�w���5��}��B���y��Ţ�Fnź	P6���:l��,����-l��e��+׵�d\v��s�#%�ދ�����nj��LH�1�?$J�Z�s�n����l��;�4~���;A����z��,�<(�9�i�X_�~��[��"�zC�����;�|�+��?�d���&��'�fb݋y�����۾�F!�9�崪�;S��O�̧��,h�V��S�t���z/~�a��L�Ɲ���S����c��2gF�����Sq�`�E�tF �B�
/Sq���O�̧��,h�V�|��-q�ٜɮpƆ�H����4H�W������������z��,S��l�ǈ�J�_�Ǉg[���ȉ�k�־/RP�C��(�l/u���!�P���sA�el$gS��:���K�ne�rE�*o.:���p�+~����f�[ۻƆeu��<̮Z;��1��h/��8��Sg3�@�<�/��NO�l����m�=�er߮��h���_�!��ZB��e�s���񱽽&O�c����)�f}Q��L�.�$��C�%tJ\a~!_�㹘eB_���]�B��Z1\3�dS����c��2gF�����XH�0�d���p�X|[��s�[~���$�M)H:aﭸ�2�������[lo�k�b�$�y�]�qs-������g%��ό�;�LȫԷ�/9�GKP�2�����Vc2�����Vcl��w&� 	���#�|"ap�� s;���*5���(ZH4~��2�����Vc2�����Vcv�iL�DH
0c`�h 1s���w�⽒���i5fqq�)/s#?�d���&�D�;E��X�\�F>>
	~�Od���E}�T��6%�6�т�H���� N��r*X]H�=7q��z��x���d��-��!1�ng�]2�nmR�#���T���I/��\]��Bjt4"�Z�X���嫋�T�%][��"��dr���L��A���)����|�Y,4�ߪ��*�/���P?Bð��T�K:+>����b~*��s�j8x��l+�Y��$|5��Җ
'x{^4��*m��L�ΪA���e�I��)G�J�cbp��'Ӡ߳A��A?�1ʤFBq��##�'�����n
V~$�x�F,*VR�U���n��뾦��q�)]Q�x��r_��m\蠓Z=�L���3f;[���p�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�o|k�Lb�5ߧE4��\�ܢ��,	սL��$����,�ǰ{�'��>b��Ќ�d2�����Vc2�����Vc�cRq>h$i�ߪOK�S]�!�I�Q�e_�UN�1�� ��2�����Vc2�����Vc����?E�p��K"]�G�D�,\ަ�It*���1��U��\�7��!��ZBk�eT�dS2O>����<��Ǉg[���Ța��k���[
�}3��*���1���Bo���+��d��Vy��h���_�!��ZB��e�s������;є:?I���\*Ծ?��CG��A:^�<���.�4�BB�U���~�*��(O"Xj�#7�E��ԛ4)�w���p���:z��j����!��ZB���E}�T�fs�歇!Ó�[���2�����Vc2�����Vc2�����Vc����'Ҥ���6��|�!7�8e�p���[�,�B2�����Vc2�����Vc2�����Vc�b+i�u�.����	�/�*�>��"������;��|B"m�ƧOAlhB" ��PK7͍��|��W&":�k�Lķ�{ �t`
�IC�oH��;��|B��EǄ���4B'�>[ӻ�ߦآ��A
�7�$G�%/���h_��s�֙L�>���+/�(�C �%;��E��٧�\�T�q�>�YŇ=�er߮�29a���Q��nj��Lk��k���d. 8��G��"�� ψ�Z;��1еQ�r�0�!7y�x�}�0�.�,E��6����|.��,�<(�9�i�X_�~��[��"�zC��s
����<����V-�łƽ�f 6j ECYz��bz���kI1C���l�q�}qj5[�*��(O"Xj�#7�E��((f��g^�W+p�ѱhkt��e�O�]�"�r�'�G�abvNx-(9�@[�_zβr�}J�DW��k���F_��_�F�'���1�FXE�>3S����x�l��15�r*Iީ�l����h���X �n�A� HX��́}H}�����Q�����M:��2��K��b��!��ZB�N4���)�Jn1�9�L�����* }�v��~nQմ�u%Y�sE��I��27bB6�_^��R������C�"�Z�X��9�R?3S����"�f7��f�mSE'h���R�ޘ�g��ra�M^���ʃh���X �^�����>�򜃗��I[�^�ґS��M�����+��~���mI��- ���X�'���-�ku�5eXL�>!�`�(i3EԔ	�8�'��P��+BY��9�
:[����>n��%+x/ �H]�毼k����<SAh�Ur��d51>�����w�!�`�(i3�022��9cbp��'Ӡ߳A��Au�����l`*��F��2vHTI�q9��Ht4 ��,� 8d�q�^!�`�(i3����~j^�q�����f-��9�K�1db��^�q:���K�n̙z7��(�^� Yv�2�����Vc2�����Vc2�����Vc�cRq>h㸁��β��L?�K<D�A���5�N^�p7N�1�� ��2�����Vc2�����Vc2�����Vc����YRwe#��`��2v]�H���'�,\ަ�It*���1���]��Y�,0��������0/����}cJQo���������k����M:��2�{�+F#J-h���X ��֞�lk��2��-����h4c�%Y�sE��I������]�^0�xP�7�gI��h"r��Zjx��7~��CF�x&��Ecc�,�[`�7���c`�\�6�(���P��
��t|q�)'������O�D� h����q*�1�pi�3h���X �{Ē�����{������٥.�*Vk������1d��2�����Vc�cRq>h$i�ߪO�5���� 3l*��2�����Vc2�����Vc_ސ����Ko˛�Y��&�D�Pk-p�󫲱�=k�Rm���X]H�=7q��z��x��<���Hn
V~$:o�>W,��q9+t�}ǆQV���C�2���R�|bd�����h�e�LD����IT#�%��-M�O��~��&V���W�V&�TA�"�Z�X�ܮI�t����q�r�nُ���f�~brw�&�z<a��N� ��M�W8߸��S�Ȍ�O��Eg׺%G*A$/q=����+'u7wO�\Vv���Z��
%��@ ��0"k��3�pڝ���hQ��g�;��|B!˕)�Lp����c6�
.�L���IJ�.߰��?�?�d���&�D�;E��Ko˛�Y��^Z���r�0h�5e��5��5DP� )Y=Wƀ?N��59X �n��n������Ut�\��ܘ[��\�!���qI/��\]��a-6�Da�X6��0Iz)զޢ:�a�79�7��{��BL��E�H�p�-a�D͢fU�9�׏�����MFi��|ր���5V��	��y��CN�I\{Hd�X4��_��t���cV��=k�Rm���|��K�iE! J�$�������e�s������Ǉ@��X��WG ���g��×�K�~�X��DL\O?H�fEd�4���z��x��ݭ/�;�J��k=�c���U!��&���`Lџ��J����	rnRͥd�ϝ�,Peal2!lL"�Z�X��NA�79)u]9�#�I�-M�O��~���N3]�nh�]#.Y��yf�ꂶ$��Q����2�nmR�#}��nd�,J�1���۪	�}a�]�w%�oφ��<�6�s�{�KrǁT8n)d�Kg�6��g���/�R�Y��/i
�\ �*؊�F��4��[=��k+��������KX��ik�����`=a�^7�-M�O��~ӊ�N6O�¼�����)�!,�!�R��q45����:s����w�4�ߪ��*�/���P?Bð��T�D<��kNgQV�.%�%���+Z�x(�i��/Rh�x#�L_�(D{ͬ�y�4����U![b��+�d��,N��w�{���á?N%��@:ND����N�&9��2B�~i�?2�nmR�#�)2?в�<H�K�,g��-A�b��LG�a�p�j8x��l+���1������[RK7ji�R�^od�~�P+���hӢ&l�ꦡ�J���(��f�x����Q�寺�Q�%��9�2�L�"Gr�v��N����b���a��c��ْ+B����>�m/4@�s Oag���e��<6C¦��_�j?�N3�J�����5��gO�q�����f-#K�v]|nkظ�����or�}�!�5����04m��hF\�肬��2a�{:��so������d���aς"�4�1|�=�5m���v��_8\/Hi����s��.��^��oF��ڵ�ڣ!�֧�ǌo�9��Cј��'P���sA��$���Xq֧�ǌo�92�ݸM�0�m�F"� 4
���֧�ǌo�9��K3��S#�F�K͕[y* }�v��~k��7'��'���Xw���e�Kfx��V$�w��9�w����������S���Q�?�M����5m���v����S�\�/�D�`���Gk��w�w u����Ug�b� ��~o��Gz��%;��E�orǟD�ui�+��V����Ca����Op�ե[�*��I�$a��@�kݵIÙ=�H�C&�����}�K�
�4l�1�¯�*k(8V�m\��ҋX����@�ڗe'�X&����ap��hٳp�VU��Jp��T���/�cͨ�@4�{����]�!����s�݀�O$��=�Q�P�TD���rs�i��s�٭��[Ø�;�x\�HP@�a����U�p��
���)󵞼�b��yv���v�x���� �N�PΚ��_q���������QV�id�F�I�~'���Xw��E֡��l{7��Z鎬�����W-O4�؏�F����U(���]�(Fw�j�@�h�β�x/�\��S)K�Ǧ��Lqc%l���`�C�����1}��xSx�lޞ�ό���.���K�Q-K��N��[B�����'���Xw�j�7����^��oF�͠Z��)2�R�wX����K�Qޡ�V�G`T�c�c��'���Xwa'�<� \�҇o"R��4�)�3�]�!���1����m��ƞQ$s�j-)�YcÐﻋ-���C�M��N�ےf����[��Z#F�Sx�lޞ�ό���.���K�Qޡ�V�G`XdF���'���Xwa'�<� \�҇o"R�Ħ�}��,�]�!���1����m��ƞQ$s�ͯ6ju�i�ﻋ-���C�M��N�ےf����[�H�x:L�Sx�lޞ�ό���.���K�Q��K���[B�����'���Xw8��;�Wx��u2�/��u��b8G_�(��hFл����'�\Vov�AT��e'���b��h�U1�\@!$m�^k�ϣ�;��p���\����ٴ��{�G��ͫ������:[2.��y�5��\��0_��@$˺/t��꫕qŧo��K�O��PJ'�`q�'�]�o Oag��!ģ{v�2O�R�<�Uh�*�bh���d��f�`��X~�.H��@�H+_��͙�W��o?�`0��	y>����g1P��/�� e8�~��<����B��B�BtQ���>Ft|�J �[�/����o��	���^�2}�0x����-Or�`�B�I&���_�Z��[���H�������b�� e8�~���5��St4!=�)-�M���V�Yct(�P:��^��g��t�[9x%UOTmc���XYo�s�#��=ҢLy\^H�����4��j2 |pD� e8�~��f��Ԡ8�tF���)e���n�`�v81⸟��0���x���"� (00�K;C�d*@��t�{�h�����#M�i�}1�O���t�t�"h�Qf�h3Z6&�<�
e���4述B���]zo}'�o�ee��&�dfl0���#�����Ź��������U-n�6j�+�W� H1����hڣ���y�e� e8�~��(-��xsF�o��ǵ�ڊ�X3U�J��K}�n���?��}?�=\e��W��4�p(q�;�$�f�RҶ=hVv��_uy�k
rx=�b��xV e8�~��G$��"�֧z���>��RN#c�&ەF9#�[��ܶ������;vLď�C����h�MCTlS�q�҇o"R\-��L�=������� e8�~����gľ�W���dx�b�W(��	!nR�K��AR%jg�Em���"B�䟷3��᧋�9ܧ!K��\4�.����|s�� �S� ���L��oI�] e8�~�� ��!~�2O�R�<�Uh�*�bh���d��f�`��X~�.H��@�H+_��͙�W��o?�`0��	yޡ�V�G`���G��� e8�~��<����B��B�BtQ���>Ft|�J �[�/����o��	���^�2}�0x����-Or�`�B�I&��kWnH=	����E�]N!aZ�Y��)�}�����T��.��W�����:��/$��H�<
o'��ȅ��Ñ���al���:S=�]KW����@_Ϳ2�t%>^��F�������{Ib!��u��Gɰ���:�#��:��L5ӥ���-���f����Oo;��$t���=�����4��lC��ۺ_~�M���g$j�SX��{��ٴ��{�G��ͫ������:[ۚܖ��`�ޡ�V�G`����g�A<�SNp>�K���y�MON|�>�)5�(���{�eV���C�T��,���G��4t���@Δ�؊�"�D���al���:S=�]KW����@_Ϳ2�t%>^��F�����ӷ�$��b!��u��Gɰ���:�#��:��L5ӥ���-���f����Oo;��$t���=�^]%S���lC��ۺ_~�M���g$j�SX��{��ٴ��{�G��ͫ������:[ۚܖ��`�ޡ�V�G`l��{[
A<�SNp>�K���y�MON|�>�)5�(���{�eV���C�T��,���G��4t�o�f{��8�؊�"�D���al���:S=�]KW����@_Ϳ2�t%>^��zN~۩qMnD�B�|d�,� �m�.�����GJR K-Ժ4� ��2�����Vc2�����Vc�d�ג��� ���>��V�"��c0�(ZH4~��2�����Vc2�����Vc@\�j�pz��Y�G�u��t�B��ꚶC�j4̗��W;��"r뾃	��s�G.5
o(=?u�AH� Ow���<�${�l'����e��G����]�w9"x�g�Hz������
���U/���I't��p �b��W'WF�K�~������hZ�tH�=���7����1g��*�s�c����t�^Z���N���D<��A[�A��l��sE���y��5�36v�( �P��Hɵ�I��<����*���al��%O&��i�n>�]Xmt<`p�ַ�sA������\�a�"�����p#9����Q��rp��U��6�����m�k�r�>?�/S�����I����=�Ŏ�yڬ�>:&���f□>�D��9]�Fk^iQ�-��^�l�,tI'��Wfe�bv={݃V5+��:��<�
�d�� }�f�ɈrS��?�d���&���{#�u����pd<H����k����ɝ\�!2A�KY�`*y�-pЊ[����oAnz��֣�:�5�D��9]�Fk^iQ��a��C���iC���0�@I��)���W�w��fD��~�Y^�������+�������zȻ�"��P�h��]XT��(Ic�!��Tӧ~-K��N��4��e/�$�*W��6����󀼐7g������¸=��tF�R�|�����&�����R y�k
rx=���7K�i�}1�O���x5xz׏�����M��ܐ�}ħ9(�z�_��������HyK�Љ���� �g�?�<2<.Xۂ!'(�`2�� �g�Aص�ٿ�MY��b֤��� �g��!`,�h��[����F�����m+�O�y�k
rx=q���:�t�>4�?J�ᡁg/V�Q�B}�����4��{�R�$�V�ޡ�V�G`9<���o4�04�jf�o��=�h�*���4�}����󀼗i�}1�O�޿�Մ*�x{^4��*m��m���.�})�?^ c��{X��@7�-�8�(�h�x#�L_�h�:��p���^�����[٩���1u4��ۂ!'(�`2����xQ�n
V~$ޡ�V�G`p��ad�J����1��`���V�{�5ߧE4��ÿR�¾B���Z#F���/9�=e$�k:~�~��@�7Л�gWaU �I}��AP:Jv��}���5�b��ۡ�y�k
rx=W��k�°eG�=:����c��>��"��a>*<UB3ޡ�V�G`���d�?�-M�O��~�W��G�t;�W���[��԰$|r9���"͵J�1��� ��U�nFޡ�V�G`�댨LV�j?U
E5��5;�`������VPY&�����R y�k
rx=�<w]��i�}1�O�߸��]
�׏�����M+�6b��1`�s䮍�����h�*�C��/y;��t����a%��w�$~��A�r��@������M�s�H�x:L�۪	�}a�]�w%�oφ��<�6�JU��j5�2�����Vc2�����Vc2�����Vc�m7���eJp�-���F#3����&�,���Fu)n2�����Vc2�����Vc2�����VcBj+)���n
2Gs�t����o*Y�kf׿����q�>�YŒ#]k�Z'�������GU4�����vIh�e�����^8�9MpW~�b��Y*��e������M:��2��!�_b�Ȳd�_�My�,L��׿��H�x:L��u����t����xe��Ok=Y�����6�c��kI1C���l�q�}qj5[!����bW��Yt�#�������\~�u.7�w�ٖE;z���������K���,tI'��WK�7R�;@�ys����ӊ[
�}3��*���1���>֐�������K]˕w���Ru-��m�3818].��@s�1�H��������	����H���,>$�'f�ٵ�e�^˯ʹ��9���v�/���ml��9�r��}�����h��%��Xcbp��'輝��eN�ħƿ�9c�Ȋ;Gx�����W���5.M+S��<FΗ�͕���/v�@ l$����\#+��S�oJ�D�=軖f�G��bu
����:�V���߃�Z�>)���t���\n	Q�1r*:����f�;�0GE�=FS�)37J*u���'��Θ/�}�<��z��}�<ͧ�:|��ΥT�t:z��j�����(�
t�ژq���U�' >�`_o��_�i��]�!��	Ǹ�y85��^�	 �wa(􆿳��Qҏ��<�q㧵�0� 0*����C˴�s� Oag�qod�֓�������/2�Q�D�{p���8
�F�:S�;��_�]�!��	Ǹ�y85��^�	 �wa(􆿳���Qs����2�`V�$�j~�����]�!��	Ǹ�y85��^�	 �wa(􆿳���Qs����F����D���pϹ7NBO��Zog����~Zh$��J�,���P���+�={"��s��(�b+�Ie�3��%b�H߫��<�dҥ��r�V��	��yF��b1�Ϋ0?���m�~����@h0�Zє���m�;bi�_��s�֙g,�e� X�]�<o����uŃp[�Ps_*�GqW�w��fD�{�����Pv��z$��?��Yn��=�gw�⽒��PAiGf;��|Bh�)���g��/e�0�o�-�W�s��={"��s��Ș�-U�6�o8:4ڜ�h���_�B�+h��:�����0h�5e��l�,ڥ�$g�[]WI�q������h���_<���Hn
V~$NgbDb�imQ���1yEI/��\]��a-6�Da�w�>���(<���w�DG\O�E朦�T�\ �͜�j�i8h��(Z+�<Vo�eo���_SJ��a�if���!#���n
V~$
3{o�[��g����s�n��뾦��q�)]Q�x��r_��m��4Ч��X�/ s f;[���p�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�o|k�Lb��ܐ�}��JdT1�V��	��y,��8v�O�w����#��X�=��'/|`��N��Z���Q���Fxkx U�_@�IX0F�M��fqwJ�D���^�MHU�:=�mI�k���(���~�7�v�ԯm��I-��]��TM���K�+EC���3��5m�-m�Z�o��q3���g����\��]+�ɸ��N��rJ�+���8ߏ[b%Ɨ��Ĥ.k�����F0D�Mv!���xx(�i��/RŻ�&ǥ��4����m1�H���W�w��fD�ޢ�}@��V���F;��|BS6=t6�Tzds�D���x�.��o� %�����b<�V5+��:��u�Y�KG�!os��qb	��G��~��<�7���1R1e�����%��s�w>o;��|B�M%>Y%��Z��0`M�Ȉ�B��ׂ4��>.g��/�ciJ�~��!8�¢5�Lm�j#%�#s��D��ð��T�K:+>�)�9K�׃]��+5u-M�O��~Ӿ9�d�L��]����YZ�[��t�ð��Th�Qf��L�zZ�K}q^J=���ɛ�?өB�R���>_|g���|��|�>�N���B�:��`{���re���?p�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�o|k�Lb��ܐ�}��JdT1�V��	��y�D�0֚ѿ8��$��dE��?'mv����1R1k� �v����ڗ�
;��|B�M%>Y%��Z��0`M�Ȉ�B��ׂ4��>.g��/�ciJ�~��!8�¢5�Lm�j#%�#s��D��ð��T�K:+>�)�9K�׃]��+5u-M�O��~Ӿ9�d�L��]����YZ�[��t�ð��Th�Qf��L�zZ�K%�줝v)��ɛ�?ө�\�G����]����Y����L9ð��Th�Qf��L�zZ�K�����-t�'+����M�g�ڄ3t���=�4�04�jfrw�&�z<a�4�ڈt׏�����M\�ܢ��,	սL��$�c�����,'t����1R1�n�S3N�.�g3Z.ӿK;�#���ᘮ�UJ%`�}lʒ^3[4JoS*�$��Pp%pv�Ka�*�W�ߟR����[��O�6 $)�lj�iE�EYZ/�W���C+���}�`��Z���Q�+�Ȋ;Gx����ZB�Ruw�C?3d�9���v�/���m�+1 v�� �tùx�Zd��䖯��l����4����q��� ��׊D��D����I�Q�#��׉󾶓�p�'Ηiu��B�A�ՙ"�z���3\0ޤ�}�����&a@ۘ36�ҋX������S8��y�)xʔ��O
�_�Z)Z�n��[��{_8�Y��=�}�Vݨ���-�9%�M(��Z��]�!��H���6D�OH��QhC��ҋX����L$�����/	� <u�}S����,�<��z��}�<ͧ�:|��ΥT�tUEcqWCl��{l�f|��:2QYeƈ�c�Z�~�����&�b<X�'���Xw���e�Kfx��V$�w�6��#�כ�������S���Q=D�I�y�6Rܝ���>�YR��j]Ln��|��L�O!f�PY�{'%s�Ǹ2���_Ma�~�Ǔ8���/��6%j_�zѩ��)�"�� )CV�v��i7N�_$�5��B>a(􆿳�k��q��־����iT u���a�Cf���P'����%���yf��>^���\�}g?	��o9���#�#99�6���0h�5e��l�,ڥ�$g�[]WI�q������h���_<���Hn
V~$X�^���܆HF4�=�I/��\]��a-6�Da9K�|���4�����g�d��%�z�J��$l���󫹬�|��{����jь$q�=�^Ey-A��{i���xȀ��D�[b%Ɨ���T��֦2��~�-�����1���#P�j2E�?�5ߧE4��c�}���Fo|k�Lbx(�i��/RŻ�&ǥ��4����m1�H���W�w��fDK�*֏�g�wj/@�'x�.��ڪ�Of���P'��NL<�E���yf��>^���\�}g?	��o9���#�#99�6���0h�5e��l�,ڥ�$g�[]WI�q������h���_<���Hn
V~$X�^���܆HF4�=�I/��\]��a-6�Da9K�|���4�����g�d��%�z�J��$l�����1�u�㤤�K��b�9f�_T(�"L?���}XO-���|��S�������<j����E����G����hK�rw�&�z<a��r����5ߧE4��p�-a�D͢fU�9�$�)�vxGY���v8N6j�"Hs��Vv�vyh�� ��г����,�ǰ�p�F�E�{���@�嗆��20�O�*C� "�w:�m�@ַ�:��ӰӬ>P�2-i_e����͂�t\	T>�I	��8����W�
J�C�7p�&'?vt��eu��q�l;1�2�-j�G�ш�g�}sۥ�Gw���#勐�E�5~09h�i�Nq�{5�h��%��Xcbp��'����Q4KҲ��r�D� �m�'�t�חEʭ�3�Jl��'p�@�JvW������(a�&�<��˰���z+/�c�Z�J
_䆼�\�v�)��+�}�+�����Ur����+��JHn��z�'>ftۿ/�>��!�F���P�sςB	5U/��@DB���h��{l�f|��rs�i�H���N���Wǖg3ȓ8���/�l|�*"k���(ӈ��";B��_�MԲ����!n}y���q���U�o=�x���Ig`i�ҋX����@�ڗe'�n�<���v�~������]�!����͙IS��⿣:�d��{l�f|�ό���.�wZ K�Ϋ�v�~������]�!��E��}����B�ip��{l�f|�ό���.�r�3P���WT�j
�I��w��,2�r@ڸWM�fx�����,@(k�n&���#��s��\.n����A�<�����y2{������Ћ�l�TUn��y{�;ۂ��IÙ=�H<}G¬x�j����)����F?2��m �A?�-��o�w_gi�.�!�����h��\�v�d����$lTǑ}�I�!?-�1~��P��~2�0�8Wn�3�RՊ��ﻋ-�����S8����ʔ?��11�g��U-�e�Y%�����F�4��W��s�2ʎ�'n�^0o**�ХM
�
Me��@ge�T�I�Lb!��u�a}��xǘ[B�����'���Xw��E���T��!�F�!n�<��Ÿ�ﻋ-�����S8�l��`�_gi�.�!����Wy����`y�������^I��}�\E��l�Q9̄�9+��z�>�C�q)ʯ���9�ǅ�k�'��P��+BY��9���$�+���)q7p�5� %�����J_�xd��j{�+F#J-��CcO^Z}��"X��[��Q[R�7�$�[ۄ���(vPZh�_ɑM��E����$�Qu𽅊"Dh\�n):��Bo�A;h�F$�Μ��VK)q7p�5jG�P�֯�^��"�c(����<m���^�b�+* �/g�d�H�RtV�^>\8�qw��UҐ�圯}Dq�f�Wဏ�R�5��a�^h�e��0�U+�qbp@�՝� s�#���k$ �Zj���
qң�:Yf�#˻��֤A|�s�X��WG ��Wr��'ǌN��,s�Q��-����!�`�(i3�H����!��8(<�'�S�|�wYð��T�ݚ�Н�!�`�(i3�ۮt@-�L�Eh��fZ���>_�����C�����"��{���m�vG)-����$�!�`�(i3!�`�(i3>\8�qw��UҐ��M��%�p@���y��lD��Z��������d�*��يC�!�`�(i3�Ra])n#���r����!�`�(i3�0e���L�Eh����N��*ȹ���Ɔ�9�ݚ�Н�!�`�(i3$f��_Ub�F�S�1 �!�`�(i3�SENan&�����R�G��m(��a(􆿳�Εq�8!�`�(i3!�`�(i3'�u�uX]�V��!����G�f��]���Rxvtm�c�oL��֬�9�^,!�`�(i3!�`�(i3Wဏ�R�5�ɣ0C��RW�7��9ᯝ
��]s��,H/��!�`�(i3���%>�rG�E`���!�`�(i3
�:qEp'{w#/ B!�`�(i3���v��\�,�6�xFg���͖n.�v�L#�?�-�Vb� �bjn� ����k��i�qs����u*w�A!�`�(i3!�`�(i3_�CE�4qްzoǸX;�%�%;a��ҜWL�!�`�(i3
�:qEp�;�P�t�5!�`�(i3$f��_Ub�F�S�1 �HN��R��bP�63Z�t��Ě���P��U@Dφ��<�6��KD���@wp ��-��Z�U9�v���O�sؤ^dN(Ҹ��j���